library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library work;
use work.FilterTypes.all;

entity FilterMemory is
  port(mem_filters : out fir_filter_array(23 downto 0));
end entity;

architecture memery of FilterMemory is
begin 
--process
--begin
  --Filter 0
  mem_filters(0)(0) <= to_signed(-13688343,32); mem_filters(0)(1) <= to_signed(9113749,32); mem_filters(0)(2) <= to_signed(-12476196,32);
  mem_filters(0)(3) <= to_signed(4577642,32); mem_filters(0)(4) <= to_signed(-7291247,32); mem_filters(0)(5) <= to_signed(-400393,32);
  mem_filters(0)(6) <= to_signed(-3976359,32); mem_filters(0)(7) <= to_signed(-4350904,32); mem_filters(0)(8) <= to_signed(-861398,32);
  mem_filters(0)(9) <= to_signed(-6691704,32); mem_filters(0)(10) <= to_signed(-530826,32); mem_filters(0)(11) <= to_signed(-7521444,32);
  mem_filters(0)(12) <= to_signed(-1075225,32); mem_filters(0)(13) <= to_signed(-6532978,32); mem_filters(0)(14) <= to_signed(-1979162,32);
  mem_filters(0)(15) <= to_signed(-4585735,32); mem_filters(0)(16) <= to_signed(-3859062,32); mem_filters(0)(17) <= to_signed(-4651511,32);
  mem_filters(0)(18) <= to_signed(-2981776,32); mem_filters(0)(19) <= to_signed(-5173432,32); mem_filters(0)(20) <= to_signed(-580120,32);
  mem_filters(0)(21) <= to_signed(-8584695,32); mem_filters(0)(22) <= to_signed(3813778,32); mem_filters(0)(23) <= to_signed(-12354092,32);
  mem_filters(0)(24) <= to_signed(7585256,32); mem_filters(0)(25) <= to_signed(-15199789,32); mem_filters(0)(26) <= to_signed(10816978,32);
  mem_filters(0)(27) <= to_signed(-15844614,32); mem_filters(0)(28) <= to_signed(10922930,32); mem_filters(0)(29) <= to_signed(-21392576,32);
  mem_filters(0)(30) <= to_signed(-17312513,32); mem_filters(0)(31) <= to_signed(-54650390,32); mem_filters(0)(32) <= to_signed(-25668014,32);
  mem_filters(0)(33) <= to_signed(-69925128,32); mem_filters(0)(34) <= to_signed(-65182760,32); mem_filters(0)(35) <= to_signed(-63405317,32);
  mem_filters(0)(36) <= to_signed(74368593,32); mem_filters(0)(37) <= to_signed(299072199,32); mem_filters(0)(38) <= to_signed(-531048362,32);
  mem_filters(0)(39) <= to_signed(-89486095,32); mem_filters(0)(40) <= to_signed(270077465,32); mem_filters(0)(41) <= to_signed(-648924392,32);
  mem_filters(0)(42) <= to_signed(-322337945,32); mem_filters(0)(43) <= to_signed(144068731,32); mem_filters(0)(44) <= to_signed(-1085206,32);
  mem_filters(0)(45) <= to_signed(-106233351,32);
  mem_filters(0)(46) <= to_signed(-21907859,32); mem_filters(0)(47) <= to_signed(104555417,32); mem_filters(0)(48) <= to_signed(115722642,32);
  mem_filters(0)(49) <= to_signed(25455963,32); mem_filters(0)(50) <= to_signed(190743375,32); mem_filters(0)(51) <= to_signed(149334428,32);
  mem_filters(0)(52) <= to_signed(-99020205,32); mem_filters(0)(53) <= to_signed(-219605552,32); mem_filters(0)(54) <= to_signed(121775271,32);
  mem_filters(0)(55) <= to_signed(129120027,32); mem_filters(0)(56) <= to_signed(22729685,32); mem_filters(0)(57) <= to_signed(-111813520,32);
  mem_filters(0)(58) <= to_signed(-170712891,32); mem_filters(0)(59) <= to_signed(77593509,32); mem_filters(0)(60) <= to_signed(-268486,32);
  mem_filters(0)(61) <= to_signed(-41472519,32); mem_filters(0)(62) <= to_signed(-30413017,32); mem_filters(0)(63) <= to_signed(24189925,32);
  mem_filters(0)(64) <= to_signed(4671803,32); mem_filters(0)(65) <= to_signed(43844810,32); mem_filters(0)(66) <= to_signed(1898167,32);
  mem_filters(0)(67) <= to_signed(41868730,32); mem_filters(0)(68) <= to_signed(65935104,32); mem_filters(0)(69) <= to_signed(16625482,32);
  mem_filters(0)(70) <= to_signed(-20738349,32); mem_filters(0)(71) <= to_signed(50171017,32); mem_filters(0)(72) <= to_signed(-3972170,32);
  mem_filters(0)(73) <= to_signed(2268576,32); mem_filters(0)(74) <= to_signed(-8039014,32); mem_filters(0)(75) <= to_signed(25904445,32);
  mem_filters(0)(76) <= to_signed(-15479535,32); mem_filters(0)(77) <= to_signed(3600221,32); mem_filters(0)(78) <= to_signed(-24958862,32);
  mem_filters(0)(79) <= to_signed(29183157,32); mem_filters(0)(80) <= to_signed(12388770,32); mem_filters(0)(81) <= to_signed(9532319,32);
  mem_filters(0)(82) <= to_signed(-4437230,32); mem_filters(0)(83) <= to_signed(-1417263,32); mem_filters(0)(84) <= to_signed(15758553,32);
  mem_filters(0)(85) <= to_signed(-2980105,32); mem_filters(0)(86) <= to_signed(1056785,32); mem_filters(0)(87) <= to_signed(-20188386,32);
  mem_filters(0)(88) <= to_signed(12228195,32); mem_filters(0)(89) <= to_signed(-10706030,32); mem_filters(0)(90) <= to_signed(8395409,32);
  mem_filters(0)(91) <= to_signed(-9498953,32); mem_filters(0)(92) <= to_signed(23027993,32); mem_filters(0)(93) <= to_signed(-9336219,32);
  mem_filters(0)(94) <= to_signed(3666831,32); mem_filters(0)(95) <= to_signed(-37629003,32); mem_filters(0)(96) <= to_signed(5453160,32);
  mem_filters(0)(97) <= to_signed(-27752691,32); mem_filters(0)(98) <= to_signed(12003648,32); mem_filters(0)(99) <= to_signed(-9003851,32);
  mem_filters(0)(100) <= to_signed(34954958,32); mem_filters(0)(101) <= to_signed(4397860,32); mem_filters(0)(102) <= to_signed(7908040,32);
  mem_filters(0)(103) <= to_signed(6073820,32); mem_filters(0)(104) <= to_signed(42573804,32); mem_filters(0)(105) <= to_signed(6379432,32);
  mem_filters(0)(106) <= to_signed(13874735,32); mem_filters(0)(107) <= to_signed(57080,32); mem_filters(0)(108) <= to_signed(-12404924,32);
  mem_filters(0)(109) <= to_signed(3972154,32); mem_filters(0)(110) <= to_signed(4466014,32); mem_filters(0)(111) <= to_signed(16054744,32);
  mem_filters(0)(112) <= to_signed(16697310,32); mem_filters(0)(113) <= to_signed(20680582,32); mem_filters(0)(114) <= to_signed(15175413,32);
  mem_filters(0)(115) <= to_signed(26836970,32); mem_filters(0)(116) <= to_signed(17308354,32); mem_filters(0)(117) <= to_signed(13252649,32);
  mem_filters(0)(118) <= to_signed(9519175,32); mem_filters(0)(119) <= to_signed(19074545,32); mem_filters(0)(120) <= to_signed(11228710,32);
  mem_filters(0)(121) <= to_signed(8532964,32); mem_filters(0)(122) <= to_signed(-2047405,32); mem_filters(0)(123) <= to_signed(4432387,32);
  mem_filters(0)(124) <= to_signed(1635373,32); mem_filters(0)(125) <= to_signed(9410221,32); mem_filters(0)(126) <= to_signed(7270717,32);
  mem_filters(0)(127) <= to_signed(5387665,32); mem_filters(0)(128) <= to_signed(2011162,32); mem_filters(0)(129) <= to_signed(3843538,32);
  mem_filters(0)(130) <= to_signed(8026176,32); mem_filters(0)(131) <= to_signed(10862632,32); mem_filters(0)(132) <= to_signed(2711394,32);
  mem_filters(0)(133) <= to_signed(4162123,32); mem_filters(0)(134) <= to_signed(-2138608,32); mem_filters(0)(135) <= to_signed(6445509,32);
  mem_filters(0)(136) <= to_signed(7298983,32); mem_filters(0)(137) <= to_signed(2488954,32); mem_filters(0)(138) <= to_signed(4699192,32);
  mem_filters(0)(139) <= to_signed(-334901,32); mem_filters(0)(140) <= to_signed(9055154,32); mem_filters(0)(141) <= to_signed(-2519086,32);
  mem_filters(0)(142) <= to_signed(10558800,32); mem_filters(0)(143) <= to_signed(795541,32); mem_filters(0)(144) <= to_signed(6729054,32);
  mem_filters(0)(145) <= to_signed(-6261900,32); mem_filters(0)(146) <= to_signed(6321185,32); mem_filters(0)(147) <= to_signed(-4381479,32);
  mem_filters(0)(148) <= to_signed(3478865,32); mem_filters(0)(149) <= to_signed(-1121564,32); mem_filters(0)(150) <= to_signed(3946110,32);
  mem_filters(0)(151) <= to_signed(-1851185,32); mem_filters(0)(152) <= to_signed(1468193,32); mem_filters(0)(153) <= to_signed(-228315,32);
  mem_filters(0)(154) <= to_signed(4409792,32); mem_filters(0)(155) <= to_signed(-1176522,32); mem_filters(0)(156) <= to_signed(2696010,32);
  mem_filters(0)(157) <= to_signed(-1707003,32); mem_filters(0)(158) <= to_signed(3114802,32); mem_filters(0)(159) <= to_signed(-2206651,32);
  mem_filters(0)(160) <= to_signed(3408097,32); mem_filters(0)(161) <= to_signed(314615,32); mem_filters(0)(162) <= to_signed(2872028,32);
  mem_filters(0)(163) <= to_signed(-1255307,32); mem_filters(0)(164) <= to_signed(-1564172,32); mem_filters(0)(165) <= to_signed(-1615050,32);
  mem_filters(0)(166) <= to_signed(-4826073,32); mem_filters(0)(167) <= to_signed(843468,32); mem_filters(0)(168) <= to_signed(-5029421,32);
  mem_filters(0)(169) <= to_signed(1787600,32); mem_filters(0)(170) <= to_signed(-8251813,32); mem_filters(0)(171) <= to_signed(1902357,32);
  mem_filters(0)(172) <= to_signed(-5560556,32); mem_filters(0)(173) <= to_signed(5079056,32); mem_filters(0)(174) <= to_signed(-5868146,32);
  mem_filters(0)(175) <= to_signed(4476898,32); mem_filters(0)(176) <= to_signed(-4537550,32); mem_filters(0)(177) <= to_signed(6744888,32);
  mem_filters(0)(178) <= to_signed(-6691636,32); mem_filters(0)(179) <= to_signed(7149877,32); mem_filters(0)(180) <= to_signed(-4498611,32);
  mem_filters(0)(181) <= to_signed(5964600,32); mem_filters(0)(182) <= to_signed(-5723303,32); mem_filters(0)(183) <= to_signed(4258156,32);
  mem_filters(0)(184) <= to_signed(-5240701,32); mem_filters(0)(185) <= to_signed(3556352,32); mem_filters(0)(186) <= to_signed(-5593858,32);
  mem_filters(0)(187) <= to_signed(7718967,32); mem_filters(0)(188) <= to_signed(-9382194,32); mem_filters(0)(189) <= to_signed(5240045,32);
  mem_filters(0)(190) <= to_signed(-10128514,32); mem_filters(0)(191) <= to_signed(10011803,32); mem_filters(0)(192) <= to_signed(-10513798,32);
  mem_filters(0)(193) <= to_signed(7597617,32); mem_filters(0)(194) <= to_signed(-12555576,32); mem_filters(0)(195) <= to_signed(10991583,32);
  mem_filters(0)(196) <= to_signed(-15508959,32); mem_filters(0)(197) <= to_signed(9439723,32); mem_filters(0)(198) <= to_signed(-16586076,32);
  mem_filters(0)(199) <= to_signed(13236605,32); mem_filters(0)(200) <= to_signed(-17875687,32); mem_filters(0)(201) <= to_signed(11533419,32);
  mem_filters(0)(202) <= to_signed(-15057789,32); mem_filters(0)(203) <= to_signed(14070081,32); mem_filters(0)(204) <= to_signed(-15656243,32);
  mem_filters(0)(205) <= to_signed(14550981,32); mem_filters(0)(206) <= to_signed(-12686020,32); mem_filters(0)(207) <= to_signed(11711278,32);
  mem_filters(0)(208) <= to_signed(-12852063,32); mem_filters(0)(209) <= to_signed(9103944,32); mem_filters(0)(210) <= to_signed(-12406565,32);
  mem_filters(0)(211) <= to_signed(5096981,32); mem_filters(0)(212) <= to_signed(-12824487,32); mem_filters(0)(213) <= to_signed(8179681,32);
  mem_filters(0)(214) <= to_signed(-7563778,32); mem_filters(0)(215) <= to_signed(3858451,32); mem_filters(0)(216) <= to_signed(-8796245,32);
  mem_filters(0)(217) <= to_signed(3181316,32); mem_filters(0)(218) <= to_signed(-4916245,32); mem_filters(0)(219) <= to_signed(219089,32);
  mem_filters(0)(220) <= to_signed(-4015410,32); mem_filters(0)(221) <= to_signed(-4480033,32); mem_filters(0)(222) <= to_signed(155240,32);
  mem_filters(0)(223) <= to_signed(-4607988,32); mem_filters(0)(224) <= to_signed(6514777,32); mem_filters(0)(225) <= to_signed(-2796003,32);
  mem_filters(0)(226) <= to_signed(10500713,32); mem_filters(0)(227) <= to_signed(-3238471,32); mem_filters(0)(228) <= to_signed(11928553,32);
  mem_filters(0)(229) <= to_signed(-11552964,32); mem_filters(0)(230) <= to_signed(3093587,32); mem_filters(0)(231) <= to_signed(-12935090,32);
  mem_filters(0)(232) <= to_signed(12613522,32); mem_filters(0)(233) <= to_signed(-3840597,32); mem_filters(0)(234) <= to_signed(8031795,32);
  mem_filters(0)(235) <= to_signed(-12521287,32); mem_filters(0)(236) <= to_signed(2125295,32); mem_filters(0)(237) <= to_signed(-13527224,32);
  mem_filters(0)(238) <= to_signed(3101573,32); mem_filters(0)(239) <= to_signed(-6388419,32); mem_filters(0)(240) <= to_signed(5717332,32);
  mem_filters(0)(241) <= to_signed(-11591945,32); mem_filters(0)(242) <= to_signed(886615,32); mem_filters(0)(243) <= to_signed(-9496735,32);
  mem_filters(0)(244) <= to_signed(7141765,32); mem_filters(0)(245) <= to_signed(-7657171,32); mem_filters(0)(246) <= to_signed(4303225,32);
  mem_filters(0)(247) <= to_signed(-5299990,32); mem_filters(0)(248) <= to_signed(-176917,32); mem_filters(0)(249) <= to_signed(-5098274,32);
  mem_filters(0)(250) <= to_signed(3071266,32); mem_filters(0)(251) <= to_signed(5458261,32); mem_filters(0)(252) <= to_signed(-396583,32);
  mem_filters(0)(253) <= to_signed(-3430368,32); mem_filters(0)(254) <= to_signed(-1825425,32); mem_filters(0)(255) <= to_signed(4774478,32);
  
  --Filter 1
  mem_filters(1)(0) <= to_signed(-7679606,32); mem_filters(1)(1) <= to_signed(3095816,32); mem_filters(1)(2) <= to_signed(-11342558,32);
  mem_filters(1)(3) <= to_signed(3681733,32); mem_filters(1)(4) <= to_signed(-12075929,32); mem_filters(1)(5) <= to_signed(2079767,32);
  mem_filters(1)(6) <= to_signed(-8787074,32); mem_filters(1)(7) <= to_signed(639277,32); mem_filters(1)(8) <= to_signed(-5496581,32);
  mem_filters(1)(9) <= to_signed(-1877398,32); mem_filters(1)(10) <= to_signed(-5903816,32); mem_filters(1)(11) <= to_signed(289825,32);
  mem_filters(1)(12) <= to_signed(-7818625,32); mem_filters(1)(13) <= to_signed(1323712,32); mem_filters(1)(14) <= to_signed(-10980032,32);
  mem_filters(1)(15) <= to_signed(4703758,32); mem_filters(1)(16) <= to_signed(-12682679,32); mem_filters(1)(17) <= to_signed(5999886,32);
  mem_filters(1)(18) <= to_signed(-15248597,32); mem_filters(1)(19) <= to_signed(9486789,32); mem_filters(1)(20) <= to_signed(-15711458,32);
  mem_filters(1)(21) <= to_signed(10288515,32); mem_filters(1)(22) <= to_signed(-15654964,32); mem_filters(1)(23) <= to_signed(11852971,32);
  mem_filters(1)(24) <= to_signed(-16173353,32); mem_filters(1)(25) <= to_signed(12773275,32); mem_filters(1)(26) <= to_signed(-28894546,32);
  mem_filters(1)(27) <= to_signed(-28371965,32); mem_filters(1)(28) <= to_signed(-72859032,32); mem_filters(1)(29) <= to_signed(-21969691,32);
  mem_filters(1)(30) <= to_signed(-109856142,32); mem_filters(1)(31) <= to_signed(-47324703,32); mem_filters(1)(32) <= to_signed(-91134528,32);
  mem_filters(1)(33) <= to_signed(239289243,32); mem_filters(1)(34) <= to_signed(266054349,32); mem_filters(1)(35) <= to_signed(-894596805,32);
  mem_filters(1)(36) <= to_signed(304690427,32); mem_filters(1)(37) <= to_signed(4103656,32); mem_filters(1)(38) <= to_signed(-948498551,32);
  mem_filters(1)(39) <= to_signed(-1291696,32); mem_filters(1)(40) <= to_signed(178921087,32); mem_filters(1)(41) <= to_signed(-37894891,32);
  mem_filters(1)(42) <= to_signed(-185275550,32); mem_filters(1)(43) <= to_signed(47775400,32); mem_filters(1)(44) <= to_signed(264987057,32);
  mem_filters(1)(45) <= to_signed(264987057,32);
  mem_filters(1)(46) <= to_signed(104857757,32); mem_filters(1)(47) <= to_signed(299515660,32); mem_filters(1)(48) <= to_signed(4526157,32);
  mem_filters(1)(49) <= to_signed(-338947622,32); mem_filters(1)(50) <= to_signed(8452720,32); mem_filters(1)(51) <= to_signed(317010592,32);
  mem_filters(1)(52) <= to_signed(26445667,32); mem_filters(1)(53) <= to_signed(-42603738,32); mem_filters(1)(54) <= to_signed(-333941577,32);
  mem_filters(1)(55) <= to_signed(130065824,32); mem_filters(1)(56) <= to_signed(62474,32); mem_filters(1)(57) <= to_signed(-10615085,32);
  mem_filters(1)(58) <= to_signed(-80263237,32); mem_filters(1)(59) <= to_signed(81254909,32); mem_filters(1)(60) <= to_signed(28203506,32);
  mem_filters(1)(61) <= to_signed(84733205,32); mem_filters(1)(62) <= to_signed(-5374172,32); mem_filters(1)(63) <= to_signed(41319589,32);
  mem_filters(1)(64) <= to_signed(78792289,32); mem_filters(1)(65) <= to_signed(-24496697,32); mem_filters(1)(66) <= to_signed(-36578382,32);
  mem_filters(1)(67) <= to_signed(78917284,32); mem_filters(1)(68) <= to_signed(23049224,32); mem_filters(1)(69) <= to_signed(-57054265,32);
  mem_filters(1)(70) <= to_signed(67897928,32); mem_filters(1)(71) <= to_signed(4846271,32); mem_filters(1)(72) <= to_signed(-17557815,32);
  mem_filters(1)(73) <= to_signed(5740257,32); mem_filters(1)(74) <= to_signed(-61327788,32); mem_filters(1)(75) <= to_signed(47010425,32);
  mem_filters(1)(76) <= to_signed(-10367325,32); mem_filters(1)(77) <= to_signed(16359795,32); mem_filters(1)(78) <= to_signed(-15467681,32);
  mem_filters(1)(79) <= to_signed(12561870,32); mem_filters(1)(80) <= to_signed(-12532625,32); mem_filters(1)(81) <= to_signed(5948617,32);
  mem_filters(1)(82) <= to_signed(-8208480,32); mem_filters(1)(83) <= to_signed(7576184,32); mem_filters(1)(84) <= to_signed(5440014,32);
  mem_filters(1)(85) <= to_signed(12185553,32); mem_filters(1)(86) <= to_signed(6144228,32); mem_filters(1)(87) <= to_signed(10710370,32);
  mem_filters(1)(88) <= to_signed(336445,32); mem_filters(1)(89) <= to_signed(20728236,32); mem_filters(1)(90) <= to_signed(-17897021,32);
  mem_filters(1)(91) <= to_signed(-11669906,32); mem_filters(1)(92) <= to_signed(-34229049,32); mem_filters(1)(93) <= to_signed(8262183,32);
  mem_filters(1)(94) <= to_signed(-10518825,32); mem_filters(1)(95) <= to_signed(37551584,32); mem_filters(1)(96) <= to_signed(24276758,32);
  mem_filters(1)(97) <= to_signed(4675992,32); mem_filters(1)(98) <= to_signed(-18135016,32); mem_filters(1)(99) <= to_signed(-2603048,32);
  mem_filters(1)(100) <= to_signed(8277585,32); mem_filters(1)(101) <= to_signed(-7085939,32); mem_filters(1)(102) <= to_signed(-406915,32);
  mem_filters(1)(103) <= to_signed(3275004,32); mem_filters(1)(104) <= to_signed(12420868,32); mem_filters(1)(105) <= to_signed(18503428,32);
  mem_filters(1)(106) <= to_signed(32114701,32); mem_filters(1)(107) <= to_signed(33528942,32); mem_filters(1)(108) <= to_signed(32761479,32);
  mem_filters(1)(109) <= to_signed(29727614,32); mem_filters(1)(110) <= to_signed(18148817,32); mem_filters(1)(111) <= to_signed(4211564,32);
  mem_filters(1)(112) <= to_signed(7351282,32); mem_filters(1)(113) <= to_signed(10869118,32); mem_filters(1)(114) <= to_signed(18996005,32);
  mem_filters(1)(115) <= to_signed(-4145825,32); mem_filters(1)(116) <= to_signed(-8127795,32); mem_filters(1)(117) <= to_signed(-11419318,32);
  mem_filters(1)(118) <= to_signed(-5547883,32); mem_filters(1)(119) <= to_signed(-1976816,32); mem_filters(1)(120) <= to_signed(2455477,32);
  mem_filters(1)(121) <= to_signed(-538421,32); mem_filters(1)(122) <= to_signed(-1980388,32); mem_filters(1)(123) <= to_signed(-3800836,32);
  mem_filters(1)(124) <= to_signed(16313801,32); mem_filters(1)(125) <= to_signed(5388146,32); mem_filters(1)(126) <= to_signed(16965945,32);
  mem_filters(1)(127) <= to_signed(1362781,32); mem_filters(1)(128) <= to_signed(16604366,32); mem_filters(1)(129) <= to_signed(4014673,32);
  mem_filters(1)(130) <= to_signed(5744945,32); mem_filters(1)(131) <= to_signed(11139638,32); mem_filters(1)(132) <= to_signed(9742538,32);
  mem_filters(1)(133) <= to_signed(9441863,32); mem_filters(1)(134) <= to_signed(-769769,32); mem_filters(1)(135) <= to_signed(10605514,32);
  mem_filters(1)(136) <= to_signed(5917564,32); mem_filters(1)(137) <= to_signed(1339303,32); mem_filters(1)(138) <= to_signed(6990763,32);
  mem_filters(1)(139) <= to_signed(4521871,32); mem_filters(1)(140) <= to_signed(14163691,32); mem_filters(1)(141) <= to_signed(-5778523,32);
  mem_filters(1)(142) <= to_signed(17204351,32); mem_filters(1)(143) <= to_signed(-2076783,32); mem_filters(1)(144) <= to_signed(13386675,32);
  mem_filters(1)(145) <= to_signed(-9625104,32); mem_filters(1)(146) <= to_signed(13971351,32); mem_filters(1)(147) <= to_signed(-2674870,32);
  mem_filters(1)(148) <= to_signed(4737901,32); mem_filters(1)(149) <= to_signed(-5603125,32); mem_filters(1)(150) <= to_signed(4322856,32);
  mem_filters(1)(151) <= to_signed(-4287512,32); mem_filters(1)(152) <= to_signed(-300028,32); mem_filters(1)(153) <= to_signed(-7000334,32);
  mem_filters(1)(154) <= to_signed(3403613,32); mem_filters(1)(155) <= to_signed(-4822288,32); mem_filters(1)(156) <= to_signed(4073617,32);
  mem_filters(1)(157) <= to_signed(-7462470,32); mem_filters(1)(158) <= to_signed(3932012,32); mem_filters(1)(159) <= to_signed(-7357260,32);
  mem_filters(1)(160) <= to_signed(5659830,32); mem_filters(1)(161) <= to_signed(-4815668,32); mem_filters(1)(162) <= to_signed(3386032,32);
  mem_filters(1)(163) <= to_signed(-5191089,32); mem_filters(1)(164) <= to_signed(2782367,32); mem_filters(1)(165) <= to_signed(1171021,32);
  mem_filters(1)(166) <= to_signed(3419674,32); mem_filters(1)(167) <= to_signed(912093,32); mem_filters(1)(168) <= to_signed(1581136,32);
  mem_filters(1)(169) <= to_signed(1024279,32); mem_filters(1)(170) <= to_signed(-59466,32); mem_filters(1)(171) <= to_signed(-1183068,32);
  mem_filters(1)(172) <= to_signed(-1043665,32); mem_filters(1)(173) <= to_signed(1978258,32); mem_filters(1)(174) <= to_signed(-3704368,32);
  mem_filters(1)(175) <= to_signed(3009743,32); mem_filters(1)(176) <= to_signed(-4218505,32); mem_filters(1)(177) <= to_signed(4140344,32);
  mem_filters(1)(178) <= to_signed(-5046171,32); mem_filters(1)(179) <= to_signed(3660782,32); mem_filters(1)(180) <= to_signed(-2103227,32);
  mem_filters(1)(181) <= to_signed(1620470,32); mem_filters(1)(182) <= to_signed(-6670241,32); mem_filters(1)(183) <= to_signed(2691128,32);
  mem_filters(1)(184) <= to_signed(-3581338,32); mem_filters(1)(185) <= to_signed(2755662,32); mem_filters(1)(186) <= to_signed(-7972747,32);
  mem_filters(1)(187) <= to_signed(3884980,32); mem_filters(1)(188) <= to_signed(-7522135,32); mem_filters(1)(189) <= to_signed(2926130,32);
  mem_filters(1)(190) <= to_signed(-11222673,32); mem_filters(1)(191) <= to_signed(6813879,32); mem_filters(1)(192) <= to_signed(-10617570,32);
  mem_filters(1)(193) <= to_signed(6456095,32); mem_filters(1)(194) <= to_signed(-11925134,32); mem_filters(1)(195) <= to_signed(5556312,32);
  mem_filters(1)(196) <= to_signed(-8457991,32); mem_filters(1)(197) <= to_signed(2011291,32); mem_filters(1)(198) <= to_signed(-7436763,32);
  mem_filters(1)(199) <= to_signed(-704976,32); mem_filters(1)(200) <= to_signed(-5730971,32); mem_filters(1)(201) <= to_signed(-2845647,32);
  mem_filters(1)(202) <= to_signed(-711136,32); mem_filters(1)(203) <= to_signed(-1811757,32); mem_filters(1)(204) <= to_signed(-2001432,32);
  mem_filters(1)(205) <= to_signed(-2861627,32); mem_filters(1)(206) <= to_signed(2972595,32); mem_filters(1)(207) <= to_signed(365130,32);
  mem_filters(1)(208) <= to_signed(-4562618,32); mem_filters(1)(209) <= to_signed(-1664814,32); mem_filters(1)(210) <= to_signed(-2858029,32);
  mem_filters(1)(211) <= to_signed(3658801,32); mem_filters(1)(212) <= to_signed(-7739861,32); mem_filters(1)(213) <= to_signed(5453437,32);
  mem_filters(1)(214) <= to_signed(-3464743,32); mem_filters(1)(215) <= to_signed(5921068,32); mem_filters(1)(216) <= to_signed(-5209926,32);
  mem_filters(1)(217) <= to_signed(3889901,32); mem_filters(1)(218) <= to_signed(-1863354,32); mem_filters(1)(219) <= to_signed(1114237,32);
  mem_filters(1)(220) <= to_signed(-1819399,32); mem_filters(1)(221) <= to_signed(218449,32); mem_filters(1)(222) <= to_signed(-4099059,32);
  mem_filters(1)(223) <= to_signed(-1738038,32); mem_filters(1)(224) <= to_signed(-2687742,32); mem_filters(1)(225) <= to_signed(5034902,32);
  mem_filters(1)(226) <= to_signed(-2352201,32); mem_filters(1)(227) <= to_signed(3663332,32); mem_filters(1)(228) <= to_signed(-2033096,32);
  mem_filters(1)(229) <= to_signed(8063177,32); mem_filters(1)(230) <= to_signed(-6914294,32); mem_filters(1)(231) <= to_signed(-2156333,32);
  mem_filters(1)(232) <= to_signed(-4621607,32); mem_filters(1)(233) <= to_signed(3734180,32); mem_filters(1)(234) <= to_signed(3668526,32);
  mem_filters(1)(235) <= to_signed(-1597505,32); mem_filters(1)(236) <= to_signed(4476403,32); mem_filters(1)(237) <= to_signed(-12702378,32);
  mem_filters(1)(238) <= to_signed(-686397,32); mem_filters(1)(239) <= to_signed(-14545228,32); mem_filters(1)(240) <= to_signed(9811758,32);
  mem_filters(1)(241) <= to_signed(-14604293,32); mem_filters(1)(242) <= to_signed(3334570,32); mem_filters(1)(243) <= to_signed(-15726690,32);
  mem_filters(1)(244) <= to_signed(8333501,32); mem_filters(1)(245) <= to_signed(-12297716,32); mem_filters(1)(246) <= to_signed(4401483,32);
  mem_filters(1)(247) <= to_signed(-8485483,32); mem_filters(1)(248) <= to_signed(5553497,32); mem_filters(1)(249) <= to_signed(-12249041,32);
  mem_filters(1)(250) <= to_signed(7373320,32); mem_filters(1)(251) <= to_signed(-4317740,32); mem_filters(1)(252) <= to_signed(19009518,32);
  mem_filters(1)(253) <= to_signed(-14211077,32); mem_filters(1)(254) <= to_signed(13722701,32); mem_filters(1)(255) <= to_signed(-16090237,32);
  
  --Filter 2
  mem_filters(2)(0) <= to_signed(-3600456,32); mem_filters(2)(1) <= to_signed(-6955322,32); mem_filters(2)(2) <= to_signed(-3154338,32);
  mem_filters(2)(3) <= to_signed(-7554761,32); mem_filters(2)(4) <= to_signed(-2314292,32); mem_filters(2)(5) <= to_signed(-6214795,32);
  mem_filters(2)(6) <= to_signed(-3132830,32); mem_filters(2)(7) <= to_signed(-5291474,32); mem_filters(2)(8) <= to_signed(-3311630,32);
  mem_filters(2)(9) <= to_signed(-2242812,32); mem_filters(2)(10) <= to_signed(-4394737,32); mem_filters(2)(11) <= to_signed(-2437418,32);
  mem_filters(2)(12) <= to_signed(-7850384,32); mem_filters(2)(13) <= to_signed(1087385,32); mem_filters(2)(14) <= to_signed(-8275493,32);
  mem_filters(2)(15) <= to_signed(950704,32); mem_filters(2)(16) <= to_signed(-10818703,32); mem_filters(2)(17) <= to_signed(3776678,32);
  mem_filters(2)(18) <= to_signed(-11851858,32); mem_filters(2)(19) <= to_signed(6195424,32); mem_filters(2)(20) <= to_signed(-13528889,32);
  mem_filters(2)(21) <= to_signed(9784588,32); mem_filters(2)(22) <= to_signed(-16465011,32); mem_filters(2)(23) <= to_signed(14925607,32);
  mem_filters(2)(24) <= to_signed(-45141154,32); mem_filters(2)(25) <= to_signed(-34155322,32); mem_filters(2)(26) <= to_signed(-95277213,32);
  mem_filters(2)(27) <= to_signed(-22257817,32); mem_filters(2)(28) <= to_signed(-151222655,32); mem_filters(2)(29) <= to_signed(-5369695,32);
  mem_filters(2)(30) <= to_signed(-130180680,32); mem_filters(2)(31) <= to_signed(473790799,32); mem_filters(2)(32) <= to_signed(-32984690,32);
  mem_filters(2)(33) <= to_signed(-842797765,32); mem_filters(2)(34) <= to_signed(510699769,32); mem_filters(2)(35) <= to_signed(-688779222,32);
  mem_filters(2)(36) <= to_signed(-605904844,32); mem_filters(2)(37) <= to_signed(136637356,32); mem_filters(2)(38) <= to_signed(93260258,32);
  mem_filters(2)(39) <= to_signed(-92819368,32); mem_filters(2)(40) <= to_signed(-178148703,32); mem_filters(2)(41) <= to_signed(393357583,32);
  mem_filters(2)(42) <= to_signed(121097143,32); mem_filters(2)(43) <= to_signed(-77843503,32); mem_filters(2)(44) <= to_signed(346115158,32);
  mem_filters(2)(45) <= to_signed(73672744,32);
  mem_filters(2)(46) <= to_signed(-205346367,32); mem_filters(2)(47) <= to_signed(-99437218,32); mem_filters(2)(48) <= to_signed(251522988,32);
  mem_filters(2)(49) <= to_signed(-93350133,32); mem_filters(2)(50) <= to_signed(57607889,32); mem_filters(2)(51) <= to_signed(-149530783,32);
  mem_filters(2)(52) <= to_signed(37553831,32); mem_filters(2)(53) <= to_signed(45820288,32); mem_filters(2)(54) <= to_signed(-35461382,32);
  mem_filters(2)(55) <= to_signed(-71595736,32); mem_filters(2)(56) <= to_signed(138390355,32); mem_filters(2)(57) <= to_signed(31449267,32);
  mem_filters(2)(58) <= to_signed(58508803,32); mem_filters(2)(59) <= to_signed(5990068,32); mem_filters(2)(60) <= to_signed(42001276,32);
  mem_filters(2)(61) <= to_signed(-45213416,32); mem_filters(2)(62) <= to_signed(76171520,32); mem_filters(2)(63) <= to_signed(-18370775,32);
  mem_filters(2)(64) <= to_signed(59832821,32); mem_filters(2)(65) <= to_signed(-65164297,32); mem_filters(2)(66) <= to_signed(46311467,32);
  mem_filters(2)(67) <= to_signed(-6067882,32); mem_filters(2)(68) <= to_signed(19186821,32); mem_filters(2)(69) <= to_signed(-11945003,32);
  mem_filters(2)(70) <= to_signed(29890296,32); mem_filters(2)(71) <= to_signed(-1593186,32); mem_filters(2)(72) <= to_signed(-9654155,32);
  mem_filters(2)(73) <= to_signed(1877644,32); mem_filters(2)(74) <= to_signed(-209339,32); mem_filters(2)(75) <= to_signed(21347802,32);
  mem_filters(2)(76) <= to_signed(-10565116,32); mem_filters(2)(77) <= to_signed(8425840,32); mem_filters(2)(78) <= to_signed(4205117,32);
  mem_filters(2)(79) <= to_signed(8364777,32); mem_filters(2)(80) <= to_signed(-9790170,32); mem_filters(2)(81) <= to_signed(5813932,32);
  mem_filters(2)(82) <= to_signed(-1228299,32); mem_filters(2)(83) <= to_signed(-6160513,32); mem_filters(2)(84) <= to_signed(413920,32);
  mem_filters(2)(85) <= to_signed(21562891,32); mem_filters(2)(86) <= to_signed(709475,32); mem_filters(2)(87) <= to_signed(-6507789,32);
  mem_filters(2)(88) <= to_signed(-2689096,32); mem_filters(2)(89) <= to_signed(470539,32); mem_filters(2)(90) <= to_signed(-6158697,32);
  mem_filters(2)(91) <= to_signed(4132398,32); mem_filters(2)(92) <= to_signed(9982775,32); mem_filters(2)(93) <= to_signed(27156462,32);
  mem_filters(2)(94) <= to_signed(12589700,32); mem_filters(2)(95) <= to_signed(-9726758,32); mem_filters(2)(96) <= to_signed(-2168170,32);
  mem_filters(2)(97) <= to_signed(2823905,32); mem_filters(2)(98) <= to_signed(-2733675,32); mem_filters(2)(99) <= to_signed(-18732836,32);
  mem_filters(2)(100) <= to_signed(4622856,32); mem_filters(2)(101) <= to_signed(6723736,32); mem_filters(2)(102) <= to_signed(18732665,32);
  mem_filters(2)(103) <= to_signed(14511796,32); mem_filters(2)(104) <= to_signed(14584395,32); mem_filters(2)(105) <= to_signed(21314636,32);
  mem_filters(2)(106) <= to_signed(24208702,32); mem_filters(2)(107) <= to_signed(16577499,32); mem_filters(2)(108) <= to_signed(998727,32);
  mem_filters(2)(109) <= to_signed(11810300,32); mem_filters(2)(110) <= to_signed(2081893,32); mem_filters(2)(111) <= to_signed(14021703,32);
  mem_filters(2)(112) <= to_signed(5988553,32); mem_filters(2)(113) <= to_signed(14927908,32); mem_filters(2)(114) <= to_signed(-2929649,32);
  mem_filters(2)(115) <= to_signed(12829232,32); mem_filters(2)(116) <= to_signed(2780174,32); mem_filters(2)(117) <= to_signed(11030709,32);
  mem_filters(2)(118) <= to_signed(-5113279,32); mem_filters(2)(119) <= to_signed(8199940,32); mem_filters(2)(120) <= to_signed(-850695,32);
  mem_filters(2)(121) <= to_signed(9477619,32); mem_filters(2)(122) <= to_signed(-1231400,32); mem_filters(2)(123) <= to_signed(2261945,32);
  mem_filters(2)(124) <= to_signed(-5296785,32); mem_filters(2)(125) <= to_signed(8599737,32); mem_filters(2)(126) <= to_signed(2932966,32);
  mem_filters(2)(127) <= to_signed(4415354,32); mem_filters(2)(128) <= to_signed(-6982220,32); mem_filters(2)(129) <= to_signed(7709870,32);
  mem_filters(2)(130) <= to_signed(2471274,32); mem_filters(2)(131) <= to_signed(11595512,32); mem_filters(2)(132) <= to_signed(-1666258,32);
  mem_filters(2)(133) <= to_signed(9316180,32); mem_filters(2)(134) <= to_signed(-4541269,32); mem_filters(2)(135) <= to_signed(18173318,32);
  mem_filters(2)(136) <= to_signed(-3150239,32); mem_filters(2)(137) <= to_signed(21999074,32); mem_filters(2)(138) <= to_signed(-7413435,32);
  mem_filters(2)(139) <= to_signed(17655288,32); mem_filters(2)(140) <= to_signed(-3972019,32); mem_filters(2)(141) <= to_signed(15222403,32);
  mem_filters(2)(142) <= to_signed(-5788641,32); mem_filters(2)(143) <= to_signed(11147595,32); mem_filters(2)(144) <= to_signed(-2640738,32);
  mem_filters(2)(145) <= to_signed(11914574,32); mem_filters(2)(146) <= to_signed(-5175827,32); mem_filters(2)(147) <= to_signed(8920667,32);
  mem_filters(2)(148) <= to_signed(-7754337,32); mem_filters(2)(149) <= to_signed(14490786,32); mem_filters(2)(150) <= to_signed(-7183749,32);
  mem_filters(2)(151) <= to_signed(12012810,32); mem_filters(2)(152) <= to_signed(-13060510,32); mem_filters(2)(153) <= to_signed(9467041,32);
  mem_filters(2)(154) <= to_signed(-8216625,32); mem_filters(2)(155) <= to_signed(9102718,32); mem_filters(2)(156) <= to_signed(-3895161,32);
  mem_filters(2)(157) <= to_signed(1428355,32); mem_filters(2)(158) <= to_signed(-4504210,32); mem_filters(2)(159) <= to_signed(-346641,32);
  mem_filters(2)(160) <= to_signed(-956540,32); mem_filters(2)(161) <= to_signed(-5799792,32); mem_filters(2)(162) <= to_signed(1173070,32);
  mem_filters(2)(163) <= to_signed(-1897433,32); mem_filters(2)(164) <= to_signed(3744594,32); mem_filters(2)(165) <= to_signed(-2903425,32);
  mem_filters(2)(166) <= to_signed(3330065,32); mem_filters(2)(167) <= to_signed(3330065,32); mem_filters(2)(168) <= to_signed(998965,32);
  mem_filters(2)(169) <= to_signed(-962192,32); mem_filters(2)(170) <= to_signed(3601268,32); mem_filters(2)(171) <= to_signed(-3434649,32);
  mem_filters(2)(172) <= to_signed(-999917,32); mem_filters(2)(173) <= to_signed(-2232928,32); mem_filters(2)(174) <= to_signed(3259791,32);
  mem_filters(2)(175) <= to_signed(-2339088,32); mem_filters(2)(176) <= to_signed(523592,32); mem_filters(2)(177) <= to_signed(-142835,32);
  mem_filters(2)(178) <= to_signed(758145,32); mem_filters(2)(179) <= to_signed(1332928,32); mem_filters(2)(180) <= to_signed(-2119259,32);
  mem_filters(2)(181) <= to_signed(4020326,32); mem_filters(2)(182) <= to_signed(-4542545,32); mem_filters(2)(183) <= to_signed(1059122,32);
  mem_filters(2)(184) <= to_signed(-7241886,32); mem_filters(2)(185) <= to_signed(2720423,32); mem_filters(2)(186) <= to_signed(-7527959,32);
  mem_filters(2)(187) <= to_signed(632554,32); mem_filters(2)(188) <= to_signed(-7965044,32); mem_filters(2)(189) <= to_signed(1675405,32);
  mem_filters(2)(190) <= to_signed(-5826009,32); mem_filters(2)(191) <= to_signed(-989232,32); mem_filters(2)(192) <= to_signed(-9212813,32);
  mem_filters(2)(193) <= to_signed(-3506908,32); mem_filters(2)(194) <= to_signed(-8602114,32); mem_filters(2)(195) <= to_signed(-3969234,32);
  mem_filters(2)(196) <= to_signed(-6069120,32); mem_filters(2)(197) <= to_signed(-3918245,32); mem_filters(2)(198) <= to_signed(-6603004,32);
  mem_filters(2)(199) <= to_signed(-3066079,32); mem_filters(2)(200) <= to_signed(-978051,32); mem_filters(2)(201) <= to_signed(-1217672,32);
  mem_filters(2)(202) <= to_signed(-5085743,32); mem_filters(2)(203) <= to_signed(-5988441,32); mem_filters(2)(204) <= to_signed(-1991215,32);
  mem_filters(2)(205) <= to_signed(-4663672,32); mem_filters(2)(206) <= to_signed(1006381,32); mem_filters(2)(207) <= to_signed(-6497991,32);
  mem_filters(2)(208) <= to_signed(4620328,32); mem_filters(2)(209) <= to_signed(-12552166,32); mem_filters(2)(210) <= to_signed(6873530,32);
  mem_filters(2)(211) <= to_signed(-9769662,32); mem_filters(2)(212) <= to_signed(11439659,32); mem_filters(2)(213) <= to_signed(-12281268,32);
  mem_filters(2)(214) <= to_signed(11402794,32); mem_filters(2)(215) <= to_signed(-7521082,32); mem_filters(2)(216) <= to_signed(8365946,32);
  mem_filters(2)(217) <= to_signed(-9898559,32); mem_filters(2)(218) <= to_signed(5265187,32); mem_filters(2)(219) <= to_signed(-5884452,32);
  mem_filters(2)(220) <= to_signed(3509131,32); mem_filters(2)(221) <= to_signed(-7997445,32); mem_filters(2)(222) <= to_signed(3277831,32);
  mem_filters(2)(223) <= to_signed(-7193211,32); mem_filters(2)(224) <= to_signed(5813596,32); mem_filters(2)(225) <= to_signed(-7199495,32);
  mem_filters(2)(226) <= to_signed(11765218,32); mem_filters(2)(227) <= to_signed(-7603384,32); mem_filters(2)(228) <= to_signed(14289047,32);
  mem_filters(2)(229) <= to_signed(-7552680,32); mem_filters(2)(230) <= to_signed(18231600,32); mem_filters(2)(231) <= to_signed(-13187401,32);
  mem_filters(2)(232) <= to_signed(6089898,32); mem_filters(2)(233) <= to_signed(-18107653,32); mem_filters(2)(234) <= to_signed(11837060,32);
  mem_filters(2)(235) <= to_signed(-10694100,32); mem_filters(2)(236) <= to_signed(9172669,32); mem_filters(2)(237) <= to_signed(-16399937,32);
  mem_filters(2)(238) <= to_signed(3043932,32); mem_filters(2)(239) <= to_signed(-21892339,32); mem_filters(2)(240) <= to_signed(3754822,32);
  mem_filters(2)(241) <= to_signed(-13943546,32); mem_filters(2)(242) <= to_signed(8645313,32); mem_filters(2)(243) <= to_signed(-19500337,32);
  mem_filters(2)(244) <= to_signed(10435171,32); mem_filters(2)(245) <= to_signed(-16729457,32); mem_filters(2)(246) <= to_signed(13011510,32);
  mem_filters(2)(247) <= to_signed(-19311921,32); mem_filters(2)(248) <= to_signed(13006600,32); mem_filters(2)(249) <= to_signed(-12623351,32);
  mem_filters(2)(250) <= to_signed(8651757,32); mem_filters(2)(251) <= to_signed(-11087108,32); mem_filters(2)(252) <= to_signed(9415045,32);
  mem_filters(2)(253) <= to_signed(-983424,32); mem_filters(2)(254) <= to_signed(2837241,32); mem_filters(2)(255) <= to_signed(-2930652,32);
  
  --Filter 3
  mem_filters(3)(0) <= to_signed(4278094,32); mem_filters(3)(1) <= to_signed(-10504447,32); mem_filters(3)(2) <= to_signed(2977939,32);
  mem_filters(3)(3) <= to_signed(-9911142,32); mem_filters(3)(4) <= to_signed(2447008,32); mem_filters(3)(5) <= to_signed(-8884512,32);
  mem_filters(3)(6) <= to_signed(-1279888,32); mem_filters(3)(7) <= to_signed(-6465049,32); mem_filters(3)(8) <= to_signed(-3941592,32);
  mem_filters(3)(9) <= to_signed(-3670103,32); mem_filters(3)(10) <= to_signed(-6148280,32); mem_filters(3)(11) <= to_signed(-392671,32);
  mem_filters(3)(12) <= to_signed(-8771284,32); mem_filters(3)(13) <= to_signed(1443009,32); mem_filters(3)(14) <= to_signed(-10375172,32);
  mem_filters(3)(15) <= to_signed(4063542,32); mem_filters(3)(16) <= to_signed(-12611595,32); mem_filters(3)(17) <= to_signed(7577142,32);
  mem_filters(3)(18) <= to_signed(-15310174,32); mem_filters(3)(19) <= to_signed(11719579,32); mem_filters(3)(20) <= to_signed(-20166698,32);
  mem_filters(3)(21) <= to_signed(18489700,32); mem_filters(3)(22) <= to_signed(-42284343,32); mem_filters(3)(23) <= to_signed(-28540930,32);
  mem_filters(3)(24) <= to_signed(-107366316,32); mem_filters(3)(25) <= to_signed(-35027289,32); mem_filters(3)(26) <= to_signed(-145546612,32);
  mem_filters(3)(27) <= to_signed(-13480730,32); mem_filters(3)(28) <= to_signed(-147547569,32); mem_filters(3)(29) <= to_signed(345104536,32);
  mem_filters(3)(30) <= to_signed(270553676,32); mem_filters(3)(31) <= to_signed(-806479082,32); mem_filters(3)(32) <= to_signed(283230423,32);
  mem_filters(3)(33) <= to_signed(-822198613,32); mem_filters(3)(34) <= to_signed(-419108166,32); mem_filters(3)(35) <= to_signed(94366589,32);
  mem_filters(3)(36) <= to_signed(-98653160,32); mem_filters(3)(37) <= to_signed(-75271301,32); mem_filters(3)(38) <= to_signed(-26412822,32);
  mem_filters(3)(39) <= to_signed(571561216,32); mem_filters(3)(40) <= to_signed(-111092955,32); mem_filters(3)(41) <= to_signed(34622239,32);
  mem_filters(3)(42) <= to_signed(221035559,32); mem_filters(3)(43) <= to_signed(33127667,32); mem_filters(3)(44) <= to_signed(-83078861,32);
  mem_filters(3)(45) <= to_signed(52815700,32);
  mem_filters(3)(46) <= to_signed(3297965,32); mem_filters(3)(47) <= to_signed(-20959497,32); mem_filters(3)(48) <= to_signed(-73702582,32);
  mem_filters(3)(49) <= to_signed(-21955379,32); mem_filters(3)(50) <= to_signed(96431361,32); mem_filters(3)(51) <= to_signed(-40984053,32);
  mem_filters(3)(52) <= to_signed(-78442251,32); mem_filters(3)(53) <= to_signed(97369312,32); mem_filters(3)(54) <= to_signed(137550282,32);
  mem_filters(3)(55) <= to_signed(90369772,32); mem_filters(3)(56) <= to_signed(18808734,32); mem_filters(3)(57) <= to_signed(-37642155,32);
  mem_filters(3)(58) <= to_signed(5160821,32); mem_filters(3)(59) <= to_signed(86034513,32); mem_filters(3)(60) <= to_signed(1193640,32);
  mem_filters(3)(61) <= to_signed(-60258463,32); mem_filters(3)(62) <= to_signed(37953907,32); mem_filters(3)(63) <= to_signed(10466277,32);
  mem_filters(3)(64) <= to_signed(-6060238,32); mem_filters(3)(65) <= to_signed(-1567701,32); mem_filters(3)(66) <= to_signed(25062799,32);
  mem_filters(3)(67) <= to_signed(5281512,32); mem_filters(3)(68) <= to_signed(-9480626,32); mem_filters(3)(69) <= to_signed(-776903,32);
  mem_filters(3)(70) <= to_signed(22270566,32); mem_filters(3)(71) <= to_signed(-512042,32); mem_filters(3)(72) <= to_signed(10805714,32);
  mem_filters(3)(73) <= to_signed(14119318,32); mem_filters(3)(74) <= to_signed(17922961,32); mem_filters(3)(75) <= to_signed(16078477,32);
  mem_filters(3)(76) <= to_signed(18867355,32); mem_filters(3)(77) <= to_signed(-22401692,32); mem_filters(3)(78) <= to_signed(20393782,32);
  mem_filters(3)(79) <= to_signed(-3619323,32); mem_filters(3)(80) <= to_signed(22531598,32); mem_filters(3)(81) <= to_signed(-14363681,32);
  mem_filters(3)(82) <= to_signed(3241628,32); mem_filters(3)(83) <= to_signed(-31623143,32); mem_filters(3)(84) <= to_signed(-7662528,32);
  mem_filters(3)(85) <= to_signed(-17306619,32); mem_filters(3)(86) <= to_signed(13069236,32); mem_filters(3)(87) <= to_signed(5556834,32);
  mem_filters(3)(88) <= to_signed(17809158,32); mem_filters(3)(89) <= to_signed(11808884,32); mem_filters(3)(90) <= to_signed(16747899,32);
  mem_filters(3)(91) <= to_signed(9260311,32); mem_filters(3)(92) <= to_signed(25572764,32); mem_filters(3)(93) <= to_signed(2666497,32);
  mem_filters(3)(94) <= to_signed(6791848,32); mem_filters(3)(95) <= to_signed(3646808,32); mem_filters(3)(96) <= to_signed(5317015,32);
  mem_filters(3)(97) <= to_signed(-18908701,32); mem_filters(3)(98) <= to_signed(-2191897,32); mem_filters(3)(99) <= to_signed(-13610382,32);
  mem_filters(3)(100) <= to_signed(785231,32); mem_filters(3)(101) <= to_signed(-14337736,32); mem_filters(3)(102) <= to_signed(12910397,32);
  mem_filters(3)(103) <= to_signed(1458539,32); mem_filters(3)(104) <= to_signed(21132730,32); mem_filters(3)(105) <= to_signed(5594422,32);
  mem_filters(3)(106) <= to_signed(27305334,32); mem_filters(3)(107) <= to_signed(12900048,32); mem_filters(3)(108) <= to_signed(26604495,32);
  mem_filters(3)(109) <= to_signed(5818730,32); mem_filters(3)(110) <= to_signed(18602419,32); mem_filters(3)(111) <= to_signed(3963153,32);
  mem_filters(3)(112) <= to_signed(5190364,32); mem_filters(3)(113) <= to_signed(470079,32); mem_filters(3)(114) <= to_signed(8970787,32);
  mem_filters(3)(115) <= to_signed(-11371171,32); mem_filters(3)(116) <= to_signed(6641773,32); mem_filters(3)(117) <= to_signed(-6365577,32);
  mem_filters(3)(118) <= to_signed(13243911,32); mem_filters(3)(119) <= to_signed(2320530,32); mem_filters(3)(120) <= to_signed(17679406,32);
  mem_filters(3)(121) <= to_signed(-7823998,32); mem_filters(3)(122) <= to_signed(7117444,32); mem_filters(3)(123) <= to_signed(8592135,32);
  mem_filters(3)(124) <= to_signed(19854029,32); mem_filters(3)(125) <= to_signed(-2090473,32); mem_filters(3)(126) <= to_signed(5384726,32);
  mem_filters(3)(127) <= to_signed(5010336,32); mem_filters(3)(128) <= to_signed(11588599,32); mem_filters(3)(129) <= to_signed(8244290,32);
  mem_filters(3)(130) <= to_signed(4599903,32); mem_filters(3)(131) <= to_signed(760664,32); mem_filters(3)(132) <= to_signed(7486753,32);
  mem_filters(3)(133) <= to_signed(4465579,32); mem_filters(3)(134) <= to_signed(6465258,32); mem_filters(3)(135) <= to_signed(3263497,32);
  mem_filters(3)(136) <= to_signed(1953045,32); mem_filters(3)(137) <= to_signed(1525746,32); mem_filters(3)(138) <= to_signed(2165239,32);
  mem_filters(3)(139) <= to_signed(9166158,32); mem_filters(3)(140) <= to_signed(-3973870,32); mem_filters(3)(141) <= to_signed(2994813,32);
  mem_filters(3)(142) <= to_signed(-7440243,32); mem_filters(3)(143) <= to_signed(7143936,32); mem_filters(3)(144) <= to_signed(-3081922,32);
  mem_filters(3)(145) <= to_signed(8477128,32); mem_filters(3)(146) <= to_signed(-3582810,32); mem_filters(3)(147) <= to_signed(5098186,32);
  mem_filters(3)(148) <= to_signed(1054605,32); mem_filters(3)(149) <= to_signed(3938656,32); mem_filters(3)(150) <= to_signed(5139105,32);
  mem_filters(3)(151) <= to_signed(-1897810,32); mem_filters(3)(152) <= to_signed(5998682,32); mem_filters(3)(153) <= to_signed(-3561541,32);
  mem_filters(3)(154) <= to_signed(7196734,32); mem_filters(3)(155) <= to_signed(-3709616,32); mem_filters(3)(156) <= to_signed(5002266,32);
  mem_filters(3)(157) <= to_signed(-2781654,32); mem_filters(3)(158) <= to_signed(1580761,32); mem_filters(3)(159) <= to_signed(-772754,32);
  mem_filters(3)(160) <= to_signed(377326,32); mem_filters(3)(161) <= to_signed(1541500,32); mem_filters(3)(162) <= to_signed(-4624502,32);
  mem_filters(3)(163) <= to_signed(3579799,32); mem_filters(3)(164) <= to_signed(-2004073,32); mem_filters(3)(165) <= to_signed(4764252,32);
  mem_filters(3)(166) <= to_signed(-870193,32); mem_filters(3)(167) <= to_signed(1638993,32); mem_filters(3)(168) <= to_signed(199354,32);
  mem_filters(3)(169) <= to_signed(2638387,32); mem_filters(3)(170) <= to_signed(1688076,32); mem_filters(3)(171) <= to_signed(4038375,32);
  mem_filters(3)(172) <= to_signed(752873,32); mem_filters(3)(173) <= to_signed(2252297,32); mem_filters(3)(174) <= to_signed(-2583039,32);
  mem_filters(3)(175) <= to_signed(4277258,32); mem_filters(3)(176) <= to_signed(-4038918,32); mem_filters(3)(177) <= to_signed(4000665,32);
  mem_filters(3)(178) <= to_signed(-6575710,32); mem_filters(3)(179) <= to_signed(5871469,32); mem_filters(3)(180) <= to_signed(-8667303,32);
  mem_filters(3)(181) <= to_signed(5621954,32); mem_filters(3)(182) <= to_signed(-8766100,32); mem_filters(3)(183) <= to_signed(6441176,32);
  mem_filters(3)(184) <= to_signed(-9546612,32); mem_filters(3)(185) <= to_signed(5553688,32); mem_filters(3)(186) <= to_signed(-7304963,32);
  mem_filters(3)(187) <= to_signed(3606648,32); mem_filters(3)(188) <= to_signed(-7739818,32); mem_filters(3)(189) <= to_signed(-1561741,32);
  mem_filters(3)(190) <= to_signed(-8237654,32); mem_filters(3)(191) <= to_signed(-4136359,32); mem_filters(3)(192) <= to_signed(-4735929,32);
  mem_filters(3)(193) <= to_signed(-8762226,32); mem_filters(3)(194) <= to_signed(-2666663,32); mem_filters(3)(195) <= to_signed(-9027434,32);
  mem_filters(3)(196) <= to_signed(-1671299,32); mem_filters(3)(197) <= to_signed(-7584214,32); mem_filters(3)(198) <= to_signed(1078219,32);
  mem_filters(3)(199) <= to_signed(-10142489,32); mem_filters(3)(200) <= to_signed(118284,32); mem_filters(3)(201) <= to_signed(-8776665,32);
  mem_filters(3)(202) <= to_signed(4968953,32); mem_filters(3)(203) <= to_signed(-7609946,32); mem_filters(3)(204) <= to_signed(2159213,32);
  mem_filters(3)(205) <= to_signed(-6877841,32); mem_filters(3)(206) <= to_signed(3250690,32); mem_filters(3)(207) <= to_signed(-6633081,32);
  mem_filters(3)(208) <= to_signed(3760365,32); mem_filters(3)(209) <= to_signed(-5290458,32); mem_filters(3)(210) <= to_signed(2654744,32);
  mem_filters(3)(211) <= to_signed(-7457562,32); mem_filters(3)(212) <= to_signed(4887743,32); mem_filters(3)(213) <= to_signed(-5241623,32);
  mem_filters(3)(214) <= to_signed(3728820,32); mem_filters(3)(215) <= to_signed(-6405116,32); mem_filters(3)(216) <= to_signed(4395043,32);
  mem_filters(3)(217) <= to_signed(-5993590,32); mem_filters(3)(218) <= to_signed(4747839,32); mem_filters(3)(219) <= to_signed(-4190825,32);
  mem_filters(3)(220) <= to_signed(4978613,32); mem_filters(3)(221) <= to_signed(-5287491,32); mem_filters(3)(222) <= to_signed(3391788,32);
  mem_filters(3)(223) <= to_signed(-5586634,32); mem_filters(3)(224) <= to_signed(4015973,32); mem_filters(3)(225) <= to_signed(-5548076,32);
  mem_filters(3)(226) <= to_signed(4562704,32); mem_filters(3)(227) <= to_signed(-8565478,32); mem_filters(3)(228) <= to_signed(7625167,32);
  mem_filters(3)(229) <= to_signed(-5157449,32); mem_filters(3)(230) <= to_signed(7987572,32); mem_filters(3)(231) <= to_signed(-4142010,32);
  mem_filters(3)(232) <= to_signed(4356129,32); mem_filters(3)(233) <= to_signed(-7904928,32); mem_filters(3)(234) <= to_signed(-3041453,32);
  mem_filters(3)(235) <= to_signed(-6402951,32); mem_filters(3)(236) <= to_signed(-2728784,32); mem_filters(3)(237) <= to_signed(-2147949,32);
  mem_filters(3)(238) <= to_signed(-335639,32); mem_filters(3)(239) <= to_signed(-3312182,32); mem_filters(3)(240) <= to_signed(-5522310,32);
  mem_filters(3)(241) <= to_signed(-10566535,32); mem_filters(3)(242) <= to_signed(-144224,32); mem_filters(3)(243) <= to_signed(-19500337,32);
  mem_filters(3)(244) <= to_signed(6079771,32); mem_filters(3)(245) <= to_signed(-6371237,32); mem_filters(3)(246) <= to_signed(1613181,32);
  mem_filters(3)(247) <= to_signed(2912986,32); mem_filters(3)(248) <= to_signed(-1905877,32); mem_filters(3)(249) <= to_signed(5827484,32);
  mem_filters(3)(250) <= to_signed(8641679,32); mem_filters(3)(251) <= to_signed(-8817292,32); mem_filters(3)(252) <= to_signed(11240434,32);
  mem_filters(3)(253) <= to_signed(-5401703,32); mem_filters(3)(254) <= to_signed(6569047,32); mem_filters(3)(255) <= to_signed(-4167002,32);
  
  --Filter 4
  mem_filters(4)(0) <= to_signed(0,32); mem_filters(4)(1) <= to_signed(0,32); mem_filters(4)(2) <= to_signed(0,32);
  mem_filters(4)(3) <= to_signed(0,32); mem_filters(4)(4) <= to_signed(0,32); mem_filters(4)(5) <= to_signed(0,32);
  mem_filters(4)(6) <= to_signed(0,32); mem_filters(4)(7) <= to_signed(0,32); mem_filters(4)(8) <= to_signed(0,32);
  mem_filters(4)(9) <= to_signed(0,32); mem_filters(4)(10) <= to_signed(0,32); mem_filters(4)(11) <= to_signed(0,32);
  mem_filters(4)(12) <= to_signed(0,32); mem_filters(4)(13) <= to_signed(0,32); mem_filters(4)(14) <= to_signed(0,32);
  mem_filters(4)(15) <= to_signed(0,32); mem_filters(4)(16) <= to_signed(0,32); mem_filters(4)(17) <= to_signed(0,32);
  mem_filters(4)(18) <= to_signed(0,32); mem_filters(4)(19) <= to_signed(0,32); mem_filters(4)(20) <= to_signed(0,32);
  mem_filters(4)(21) <= to_signed(0,32); mem_filters(4)(22) <= to_signed(0,32); mem_filters(4)(23) <= to_signed(0,32);
  mem_filters(4)(24) <= to_signed(0,32); mem_filters(4)(25) <= to_signed(0,32); mem_filters(4)(26) <= to_signed(0,32);
  mem_filters(4)(27) <= to_signed(0,32); mem_filters(4)(28) <= to_signed(0,32); mem_filters(4)(29) <= to_signed(0,32);
  mem_filters(4)(30) <= to_signed(0,32); mem_filters(4)(31) <= to_signed(0,32); mem_filters(4)(32) <= to_signed(0,32);
  mem_filters(4)(33) <= to_signed(0,32); mem_filters(4)(34) <= to_signed(0,32); mem_filters(4)(35) <= to_signed(0,32);
  mem_filters(4)(36) <= to_signed(0,32); mem_filters(4)(37) <= to_signed(0,32); mem_filters(4)(38) <= to_signed(0,32);
  mem_filters(4)(39) <= to_signed(0,32); mem_filters(4)(40) <= to_signed(0,32); mem_filters(4)(41) <= to_signed(0,32);
  mem_filters(4)(42) <= to_signed(0,32); mem_filters(4)(43) <= to_signed(0,32); mem_filters(4)(44) <= to_signed(0,32);
  mem_filters(4)(45) <= to_signed(0,32);
  mem_filters(4)(46) <= to_signed(0,32); mem_filters(4)(47) <= to_signed(0,32); mem_filters(4)(48) <= to_signed(0,32);
  mem_filters(4)(49) <= to_signed(0,32); mem_filters(4)(50) <= to_signed(0,32); mem_filters(4)(51) <= to_signed(0,32);
  mem_filters(4)(52) <= to_signed(0,32); mem_filters(4)(53) <= to_signed(0,32); mem_filters(4)(54) <= to_signed(0,32);
  mem_filters(4)(55) <= to_signed(0,32); mem_filters(4)(56) <= to_signed(0,32); mem_filters(4)(57) <= to_signed(0,32);
  mem_filters(4)(58) <= to_signed(0,32); mem_filters(4)(59) <= to_signed(0,32); mem_filters(4)(60) <= to_signed(0,32);
  mem_filters(4)(61) <= to_signed(0,32); mem_filters(4)(62) <= to_signed(0,32); mem_filters(4)(63) <= to_signed(0,32);
  mem_filters(4)(64) <= to_signed(0,32); mem_filters(4)(65) <= to_signed(0,32); mem_filters(4)(66) <= to_signed(0,32);
  mem_filters(4)(67) <= to_signed(0,32); mem_filters(4)(68) <= to_signed(0,32); mem_filters(4)(69) <= to_signed(0,32);
  mem_filters(4)(70) <= to_signed(0,32); mem_filters(4)(71) <= to_signed(0,32); mem_filters(4)(72) <= to_signed(0,32);
  mem_filters(4)(73) <= to_signed(0,32); mem_filters(4)(74) <= to_signed(0,32); mem_filters(4)(75) <= to_signed(0,32);
  mem_filters(4)(76) <= to_signed(0,32); mem_filters(4)(77) <= to_signed(0,32); mem_filters(4)(78) <= to_signed(0,32);
  mem_filters(4)(79) <= to_signed(0,32); mem_filters(4)(80) <= to_signed(0,32); mem_filters(4)(81) <= to_signed(0,32);
  mem_filters(4)(82) <= to_signed(0,32); mem_filters(4)(83) <= to_signed(0,32); mem_filters(4)(84) <= to_signed(0,32);
  mem_filters(4)(85) <= to_signed(0,32); mem_filters(4)(86) <= to_signed(0,32); mem_filters(4)(87) <= to_signed(0,32);
  mem_filters(4)(88) <= to_signed(0,32); mem_filters(4)(89) <= to_signed(0,32); mem_filters(4)(90) <= to_signed(0,32);
  mem_filters(4)(91) <= to_signed(0,32); mem_filters(4)(92) <= to_signed(0,32); mem_filters(4)(93) <= to_signed(0,32);
  mem_filters(4)(94) <= to_signed(0,32); mem_filters(4)(95) <= to_signed(0,32); mem_filters(4)(96) <= to_signed(0,32);
  mem_filters(4)(97) <= to_signed(0,32); mem_filters(4)(98) <= to_signed(0,32); mem_filters(4)(99) <= to_signed(0,32);
  mem_filters(4)(100) <= to_signed(0,32); mem_filters(4)(101) <= to_signed(0,32); mem_filters(4)(102) <= to_signed(0,32);
  mem_filters(4)(103) <= to_signed(0,32); mem_filters(4)(104) <= to_signed(0,32); mem_filters(4)(105) <= to_signed(0,32);
  mem_filters(4)(106) <= to_signed(0,32); mem_filters(4)(107) <= to_signed(0,32); mem_filters(4)(108) <= to_signed(0,32);
  mem_filters(4)(109) <= to_signed(0,32); mem_filters(4)(110) <= to_signed(0,32); mem_filters(4)(111) <= to_signed(0,32);
  mem_filters(4)(112) <= to_signed(0,32); mem_filters(4)(113) <= to_signed(0,32); mem_filters(4)(114) <= to_signed(0,32);
  mem_filters(4)(115) <= to_signed(0,32); mem_filters(4)(116) <= to_signed(0,32); mem_filters(4)(117) <= to_signed(0,32);
  mem_filters(4)(118) <= to_signed(0,32); mem_filters(4)(119) <= to_signed(0,32); mem_filters(4)(120) <= to_signed(0,32);
  mem_filters(4)(121) <= to_signed(0,32); mem_filters(4)(122) <= to_signed(0,32); mem_filters(4)(123) <= to_signed(0,32);
  mem_filters(4)(124) <= to_signed(0,32); mem_filters(4)(125) <= to_signed(0,32); mem_filters(4)(126) <= to_signed(0,32);
  mem_filters(4)(127) <= to_signed(0,32); mem_filters(4)(128) <= to_signed(0,32); mem_filters(4)(129) <= to_signed(0,32);
  mem_filters(4)(130) <= to_signed(0,32); mem_filters(4)(131) <= to_signed(0,32); mem_filters(4)(132) <= to_signed(0,32);
  mem_filters(4)(133) <= to_signed(0,32); mem_filters(4)(134) <= to_signed(0,32); mem_filters(4)(135) <= to_signed(0,32);
  mem_filters(4)(136) <= to_signed(0,32); mem_filters(4)(137) <= to_signed(0,32); mem_filters(4)(138) <= to_signed(0,32);
  mem_filters(4)(139) <= to_signed(0,32); mem_filters(4)(140) <= to_signed(0,32); mem_filters(4)(141) <= to_signed(0,32);
  mem_filters(4)(142) <= to_signed(0,32); mem_filters(4)(143) <= to_signed(0,32); mem_filters(4)(144) <= to_signed(0,32);
  mem_filters(4)(145) <= to_signed(0,32); mem_filters(4)(146) <= to_signed(0,32); mem_filters(4)(147) <= to_signed(0,32);
  mem_filters(4)(148) <= to_signed(0,32); mem_filters(4)(149) <= to_signed(0,32); mem_filters(4)(150) <= to_signed(0,32);
  mem_filters(4)(151) <= to_signed(0,32); mem_filters(4)(152) <= to_signed(0,32); mem_filters(4)(153) <= to_signed(0,32);
  mem_filters(4)(154) <= to_signed(0,32); mem_filters(4)(155) <= to_signed(0,32); mem_filters(4)(156) <= to_signed(0,32);
  mem_filters(4)(157) <= to_signed(0,32); mem_filters(4)(158) <= to_signed(0,32); mem_filters(4)(159) <= to_signed(0,32);
  mem_filters(4)(160) <= to_signed(0,32); mem_filters(4)(161) <= to_signed(0,32); mem_filters(4)(162) <= to_signed(0,32);
  mem_filters(4)(163) <= to_signed(0,32); mem_filters(4)(164) <= to_signed(0,32); mem_filters(4)(165) <= to_signed(0,32);
  mem_filters(4)(166) <= to_signed(0,32); mem_filters(4)(167) <= to_signed(0,32); mem_filters(4)(168) <= to_signed(0,32);
  mem_filters(4)(169) <= to_signed(0,32); mem_filters(4)(170) <= to_signed(0,32); mem_filters(4)(171) <= to_signed(0,32);
  mem_filters(4)(172) <= to_signed(0,32); mem_filters(4)(173) <= to_signed(0,32); mem_filters(4)(174) <= to_signed(0,32);
  mem_filters(4)(175) <= to_signed(0,32); mem_filters(4)(176) <= to_signed(0,32); mem_filters(4)(177) <= to_signed(0,32);
  mem_filters(4)(178) <= to_signed(0,32); mem_filters(4)(179) <= to_signed(0,32); mem_filters(4)(180) <= to_signed(0,32);
  mem_filters(4)(181) <= to_signed(0,32); mem_filters(4)(182) <= to_signed(0,32); mem_filters(4)(183) <= to_signed(0,32);
  mem_filters(4)(184) <= to_signed(0,32); mem_filters(4)(185) <= to_signed(0,32); mem_filters(4)(186) <= to_signed(0,32);
  mem_filters(4)(187) <= to_signed(0,32); mem_filters(4)(188) <= to_signed(0,32); mem_filters(4)(189) <= to_signed(0,32);
  mem_filters(4)(190) <= to_signed(0,32); mem_filters(4)(191) <= to_signed(0,32); mem_filters(4)(192) <= to_signed(0,32);
  mem_filters(4)(193) <= to_signed(0,32); mem_filters(4)(194) <= to_signed(0,32); mem_filters(4)(195) <= to_signed(0,32);
  mem_filters(4)(196) <= to_signed(0,32); mem_filters(4)(197) <= to_signed(0,32); mem_filters(4)(198) <= to_signed(0,32);
  mem_filters(4)(199) <= to_signed(0,32); mem_filters(4)(200) <= to_signed(0,32); mem_filters(4)(201) <= to_signed(0,32);
  mem_filters(4)(202) <= to_signed(0,32); mem_filters(4)(203) <= to_signed(0,32); mem_filters(4)(204) <= to_signed(0,32);
  mem_filters(4)(205) <= to_signed(0,32); mem_filters(4)(206) <= to_signed(0,32); mem_filters(4)(207) <= to_signed(0,32);
  mem_filters(4)(208) <= to_signed(0,32); mem_filters(4)(209) <= to_signed(0,32); mem_filters(4)(210) <= to_signed(0,32);
  mem_filters(4)(211) <= to_signed(0,32); mem_filters(4)(212) <= to_signed(0,32); mem_filters(4)(213) <= to_signed(0,32);
  mem_filters(4)(214) <= to_signed(0,32); mem_filters(4)(215) <= to_signed(0,32); mem_filters(4)(216) <= to_signed(0,32);
  mem_filters(4)(217) <= to_signed(0,32); mem_filters(4)(218) <= to_signed(0,32); mem_filters(4)(219) <= to_signed(0,32);
  mem_filters(4)(220) <= to_signed(0,32); mem_filters(4)(221) <= to_signed(0,32); mem_filters(4)(222) <= to_signed(0,32);
  mem_filters(4)(223) <= to_signed(0,32); mem_filters(4)(224) <= to_signed(0,32); mem_filters(4)(225) <= to_signed(0,32);
  mem_filters(4)(226) <= to_signed(0,32); mem_filters(4)(227) <= to_signed(0,32); mem_filters(4)(228) <= to_signed(0,32);
  mem_filters(4)(229) <= to_signed(0,32); mem_filters(4)(230) <= to_signed(0,32); mem_filters(4)(231) <= to_signed(0,32);
  mem_filters(4)(232) <= to_signed(0,32); mem_filters(4)(233) <= to_signed(0,32); mem_filters(4)(234) <= to_signed(0,32);
  mem_filters(4)(235) <= to_signed(0,32); mem_filters(4)(236) <= to_signed(0,32); mem_filters(4)(237) <= to_signed(0,32);
  mem_filters(4)(238) <= to_signed(0,32); mem_filters(4)(239) <= to_signed(0,32); mem_filters(4)(240) <= to_signed(0,32);
  mem_filters(4)(241) <= to_signed(0,32); mem_filters(4)(242) <= to_signed(0,32); mem_filters(4)(243) <= to_signed(0,32);
  mem_filters(4)(244) <= to_signed(0,32); mem_filters(4)(245) <= to_signed(0,32); mem_filters(4)(246) <= to_signed(0,32);
  mem_filters(4)(247) <= to_signed(0,32); mem_filters(4)(248) <= to_signed(0,32); mem_filters(4)(249) <= to_signed(0,32);
  mem_filters(4)(250) <= to_signed(0,32); mem_filters(4)(251) <= to_signed(0,32); mem_filters(4)(252) <= to_signed(0,32);
  mem_filters(4)(253) <= to_signed(0,32); mem_filters(4)(254) <= to_signed(0,32); mem_filters(4)(255) <= to_signed(0,32);
  
  --Filter 5
  mem_filters(5)(0) <= to_signed(0,32); mem_filters(5)(1) <= to_signed(0,32); mem_filters(5)(2) <= to_signed(0,32);
  mem_filters(5)(3) <= to_signed(0,32); mem_filters(5)(4) <= to_signed(0,32); mem_filters(5)(5) <= to_signed(0,32);
  mem_filters(5)(6) <= to_signed(0,32); mem_filters(5)(7) <= to_signed(0,32); mem_filters(5)(8) <= to_signed(0,32);
  mem_filters(5)(9) <= to_signed(0,32); mem_filters(5)(10) <= to_signed(0,32); mem_filters(5)(11) <= to_signed(0,32);
  mem_filters(5)(12) <= to_signed(0,32); mem_filters(5)(13) <= to_signed(0,32); mem_filters(5)(14) <= to_signed(0,32);
  mem_filters(5)(15) <= to_signed(0,32); mem_filters(5)(16) <= to_signed(0,32); mem_filters(5)(17) <= to_signed(0,32);
  mem_filters(5)(18) <= to_signed(0,32); mem_filters(5)(19) <= to_signed(0,32); mem_filters(5)(20) <= to_signed(0,32);
  mem_filters(5)(21) <= to_signed(0,32); mem_filters(5)(22) <= to_signed(0,32); mem_filters(5)(23) <= to_signed(0,32);
  mem_filters(5)(24) <= to_signed(0,32); mem_filters(5)(25) <= to_signed(0,32); mem_filters(5)(26) <= to_signed(0,32);
  mem_filters(5)(27) <= to_signed(0,32); mem_filters(5)(28) <= to_signed(0,32); mem_filters(5)(29) <= to_signed(0,32);
  mem_filters(5)(30) <= to_signed(0,32); mem_filters(5)(31) <= to_signed(0,32); mem_filters(5)(32) <= to_signed(0,32);
  mem_filters(5)(33) <= to_signed(0,32); mem_filters(5)(34) <= to_signed(0,32); mem_filters(5)(35) <= to_signed(0,32);
  mem_filters(5)(36) <= to_signed(0,32); mem_filters(5)(37) <= to_signed(0,32); mem_filters(5)(38) <= to_signed(0,32);
  mem_filters(5)(39) <= to_signed(0,32); mem_filters(5)(40) <= to_signed(0,32); mem_filters(5)(41) <= to_signed(0,32);
  mem_filters(5)(42) <= to_signed(0,32); mem_filters(5)(43) <= to_signed(0,32); mem_filters(5)(44) <= to_signed(0,32);
  mem_filters(5)(45) <= to_signed(0,32);
  mem_filters(5)(46) <= to_signed(0,32); mem_filters(5)(47) <= to_signed(0,32); mem_filters(5)(48) <= to_signed(0,32);
  mem_filters(5)(49) <= to_signed(0,32); mem_filters(5)(50) <= to_signed(0,32); mem_filters(5)(51) <= to_signed(0,32);
  mem_filters(5)(52) <= to_signed(0,32); mem_filters(5)(53) <= to_signed(0,32); mem_filters(5)(54) <= to_signed(0,32);
  mem_filters(5)(55) <= to_signed(0,32); mem_filters(5)(56) <= to_signed(0,32); mem_filters(5)(57) <= to_signed(0,32);
  mem_filters(5)(58) <= to_signed(0,32); mem_filters(5)(59) <= to_signed(0,32); mem_filters(5)(60) <= to_signed(0,32);
  mem_filters(5)(61) <= to_signed(0,32); mem_filters(5)(62) <= to_signed(0,32); mem_filters(5)(63) <= to_signed(0,32);
  mem_filters(5)(64) <= to_signed(0,32); mem_filters(5)(65) <= to_signed(0,32); mem_filters(5)(66) <= to_signed(0,32);
  mem_filters(5)(67) <= to_signed(0,32); mem_filters(5)(68) <= to_signed(0,32); mem_filters(5)(69) <= to_signed(0,32);
  mem_filters(5)(70) <= to_signed(0,32); mem_filters(5)(71) <= to_signed(0,32); mem_filters(5)(72) <= to_signed(0,32);
  mem_filters(5)(73) <= to_signed(0,32); mem_filters(5)(74) <= to_signed(0,32); mem_filters(5)(75) <= to_signed(0,32);
  mem_filters(5)(76) <= to_signed(0,32); mem_filters(5)(77) <= to_signed(0,32); mem_filters(5)(78) <= to_signed(0,32);
  mem_filters(5)(79) <= to_signed(0,32); mem_filters(5)(80) <= to_signed(0,32); mem_filters(5)(81) <= to_signed(0,32);
  mem_filters(5)(82) <= to_signed(0,32); mem_filters(5)(83) <= to_signed(0,32); mem_filters(5)(84) <= to_signed(0,32);
  mem_filters(5)(85) <= to_signed(0,32); mem_filters(5)(86) <= to_signed(0,32); mem_filters(5)(87) <= to_signed(0,32);
  mem_filters(5)(88) <= to_signed(0,32); mem_filters(5)(89) <= to_signed(0,32); mem_filters(5)(90) <= to_signed(0,32);
  mem_filters(5)(91) <= to_signed(0,32); mem_filters(5)(92) <= to_signed(0,32); mem_filters(5)(93) <= to_signed(0,32);
  mem_filters(5)(94) <= to_signed(0,32); mem_filters(5)(95) <= to_signed(0,32); mem_filters(5)(96) <= to_signed(0,32);
  mem_filters(5)(97) <= to_signed(0,32); mem_filters(5)(98) <= to_signed(0,32); mem_filters(5)(99) <= to_signed(0,32);
  mem_filters(5)(100) <= to_signed(0,32); mem_filters(5)(101) <= to_signed(0,32); mem_filters(5)(102) <= to_signed(0,32);
  mem_filters(5)(103) <= to_signed(0,32); mem_filters(5)(104) <= to_signed(0,32); mem_filters(5)(105) <= to_signed(0,32);
  mem_filters(5)(106) <= to_signed(0,32); mem_filters(5)(107) <= to_signed(0,32); mem_filters(5)(108) <= to_signed(0,32);
  mem_filters(5)(109) <= to_signed(0,32); mem_filters(5)(110) <= to_signed(0,32); mem_filters(5)(111) <= to_signed(0,32);
  mem_filters(5)(112) <= to_signed(0,32); mem_filters(5)(113) <= to_signed(0,32); mem_filters(5)(114) <= to_signed(0,32);
  mem_filters(5)(115) <= to_signed(0,32); mem_filters(5)(116) <= to_signed(0,32); mem_filters(5)(117) <= to_signed(0,32);
  mem_filters(5)(118) <= to_signed(0,32); mem_filters(5)(119) <= to_signed(0,32); mem_filters(5)(120) <= to_signed(0,32);
  mem_filters(5)(121) <= to_signed(0,32); mem_filters(5)(122) <= to_signed(0,32); mem_filters(5)(123) <= to_signed(0,32);
  mem_filters(5)(124) <= to_signed(0,32); mem_filters(5)(125) <= to_signed(0,32); mem_filters(5)(126) <= to_signed(0,32);
  mem_filters(5)(127) <= to_signed(0,32); mem_filters(5)(128) <= to_signed(0,32); mem_filters(5)(129) <= to_signed(0,32);
  mem_filters(5)(130) <= to_signed(0,32); mem_filters(5)(131) <= to_signed(0,32); mem_filters(5)(132) <= to_signed(0,32);
  mem_filters(5)(133) <= to_signed(0,32); mem_filters(5)(134) <= to_signed(0,32); mem_filters(5)(135) <= to_signed(0,32);
  mem_filters(5)(136) <= to_signed(0,32); mem_filters(5)(137) <= to_signed(0,32); mem_filters(5)(138) <= to_signed(0,32);
  mem_filters(5)(139) <= to_signed(0,32); mem_filters(5)(140) <= to_signed(0,32); mem_filters(5)(141) <= to_signed(0,32);
  mem_filters(5)(142) <= to_signed(0,32); mem_filters(5)(143) <= to_signed(0,32); mem_filters(5)(144) <= to_signed(0,32);
  mem_filters(5)(145) <= to_signed(0,32); mem_filters(5)(146) <= to_signed(0,32); mem_filters(5)(147) <= to_signed(0,32);
  mem_filters(5)(148) <= to_signed(0,32); mem_filters(5)(149) <= to_signed(0,32); mem_filters(5)(150) <= to_signed(0,32);
  mem_filters(5)(151) <= to_signed(0,32); mem_filters(5)(152) <= to_signed(0,32); mem_filters(5)(153) <= to_signed(0,32);
  mem_filters(5)(154) <= to_signed(0,32); mem_filters(5)(155) <= to_signed(0,32); mem_filters(5)(156) <= to_signed(0,32);
  mem_filters(5)(157) <= to_signed(0,32); mem_filters(5)(158) <= to_signed(0,32); mem_filters(5)(159) <= to_signed(0,32);
  mem_filters(5)(160) <= to_signed(0,32); mem_filters(5)(161) <= to_signed(0,32); mem_filters(5)(162) <= to_signed(0,32);
  mem_filters(5)(163) <= to_signed(0,32); mem_filters(5)(164) <= to_signed(0,32); mem_filters(5)(165) <= to_signed(0,32);
  mem_filters(5)(166) <= to_signed(0,32); mem_filters(5)(167) <= to_signed(0,32); mem_filters(5)(168) <= to_signed(0,32);
  mem_filters(5)(169) <= to_signed(0,32); mem_filters(5)(170) <= to_signed(0,32); mem_filters(5)(171) <= to_signed(0,32);
  mem_filters(5)(172) <= to_signed(0,32); mem_filters(5)(173) <= to_signed(0,32); mem_filters(5)(174) <= to_signed(0,32);
  mem_filters(5)(175) <= to_signed(0,32); mem_filters(5)(176) <= to_signed(0,32); mem_filters(5)(177) <= to_signed(0,32);
  mem_filters(5)(178) <= to_signed(0,32); mem_filters(5)(179) <= to_signed(0,32); mem_filters(5)(180) <= to_signed(0,32);
  mem_filters(5)(181) <= to_signed(0,32); mem_filters(5)(182) <= to_signed(0,32); mem_filters(5)(183) <= to_signed(0,32);
  mem_filters(5)(184) <= to_signed(0,32); mem_filters(5)(185) <= to_signed(0,32); mem_filters(5)(186) <= to_signed(0,32);
  mem_filters(5)(187) <= to_signed(0,32); mem_filters(5)(188) <= to_signed(0,32); mem_filters(5)(189) <= to_signed(0,32);
  mem_filters(5)(190) <= to_signed(0,32); mem_filters(5)(191) <= to_signed(0,32); mem_filters(5)(192) <= to_signed(0,32);
  mem_filters(5)(193) <= to_signed(0,32); mem_filters(5)(194) <= to_signed(0,32); mem_filters(5)(195) <= to_signed(0,32);
  mem_filters(5)(196) <= to_signed(0,32); mem_filters(5)(197) <= to_signed(0,32); mem_filters(5)(198) <= to_signed(0,32);
  mem_filters(5)(199) <= to_signed(0,32); mem_filters(5)(200) <= to_signed(0,32); mem_filters(5)(201) <= to_signed(0,32);
  mem_filters(5)(202) <= to_signed(0,32); mem_filters(5)(203) <= to_signed(0,32); mem_filters(5)(204) <= to_signed(0,32);
  mem_filters(5)(205) <= to_signed(0,32); mem_filters(5)(206) <= to_signed(0,32); mem_filters(5)(207) <= to_signed(0,32);
  mem_filters(5)(208) <= to_signed(0,32); mem_filters(5)(209) <= to_signed(0,32); mem_filters(5)(210) <= to_signed(0,32);
  mem_filters(5)(211) <= to_signed(0,32); mem_filters(5)(212) <= to_signed(0,32); mem_filters(5)(213) <= to_signed(0,32);
  mem_filters(5)(214) <= to_signed(0,32); mem_filters(5)(215) <= to_signed(0,32); mem_filters(5)(216) <= to_signed(0,32);
  mem_filters(5)(217) <= to_signed(0,32); mem_filters(5)(218) <= to_signed(0,32); mem_filters(5)(219) <= to_signed(0,32);
  mem_filters(5)(220) <= to_signed(0,32); mem_filters(5)(221) <= to_signed(0,32); mem_filters(5)(222) <= to_signed(0,32);
  mem_filters(5)(223) <= to_signed(0,32); mem_filters(5)(224) <= to_signed(0,32); mem_filters(5)(225) <= to_signed(0,32);
  mem_filters(5)(226) <= to_signed(0,32); mem_filters(5)(227) <= to_signed(0,32); mem_filters(5)(228) <= to_signed(0,32);
  mem_filters(5)(229) <= to_signed(0,32); mem_filters(5)(230) <= to_signed(0,32); mem_filters(5)(231) <= to_signed(0,32);
  mem_filters(5)(232) <= to_signed(0,32); mem_filters(5)(233) <= to_signed(0,32); mem_filters(5)(234) <= to_signed(0,32);
  mem_filters(5)(235) <= to_signed(0,32); mem_filters(5)(236) <= to_signed(0,32); mem_filters(5)(237) <= to_signed(0,32);
  mem_filters(5)(238) <= to_signed(0,32); mem_filters(5)(239) <= to_signed(0,32); mem_filters(5)(240) <= to_signed(0,32);
  mem_filters(5)(241) <= to_signed(0,32); mem_filters(5)(242) <= to_signed(0,32); mem_filters(5)(243) <= to_signed(0,32);
  mem_filters(5)(244) <= to_signed(0,32); mem_filters(5)(245) <= to_signed(0,32); mem_filters(5)(246) <= to_signed(0,32);
  mem_filters(5)(247) <= to_signed(0,32); mem_filters(5)(248) <= to_signed(0,32); mem_filters(5)(249) <= to_signed(0,32);
  mem_filters(5)(250) <= to_signed(0,32); mem_filters(5)(251) <= to_signed(0,32); mem_filters(5)(252) <= to_signed(0,32);
  mem_filters(5)(253) <= to_signed(0,32); mem_filters(5)(254) <= to_signed(0,32); mem_filters(5)(255) <= to_signed(0,32);
  
  --Filter 6
  mem_filters(6)(0) <= to_signed(0,32); mem_filters(6)(1) <= to_signed(0,32); mem_filters(6)(2) <= to_signed(0,32);
  mem_filters(6)(3) <= to_signed(0,32); mem_filters(6)(4) <= to_signed(0,32); mem_filters(6)(5) <= to_signed(0,32);
  mem_filters(6)(6) <= to_signed(0,32); mem_filters(6)(7) <= to_signed(0,32); mem_filters(6)(8) <= to_signed(0,32);
  mem_filters(6)(9) <= to_signed(0,32); mem_filters(6)(10) <= to_signed(0,32); mem_filters(6)(11) <= to_signed(0,32);
  mem_filters(6)(12) <= to_signed(0,32); mem_filters(6)(13) <= to_signed(0,32); mem_filters(6)(14) <= to_signed(0,32);
  mem_filters(6)(15) <= to_signed(0,32); mem_filters(6)(16) <= to_signed(0,32); mem_filters(6)(17) <= to_signed(0,32);
  mem_filters(6)(18) <= to_signed(0,32); mem_filters(6)(19) <= to_signed(0,32); mem_filters(6)(20) <= to_signed(0,32);
  mem_filters(6)(21) <= to_signed(0,32); mem_filters(6)(22) <= to_signed(0,32); mem_filters(6)(23) <= to_signed(0,32);
  mem_filters(6)(24) <= to_signed(0,32); mem_filters(6)(25) <= to_signed(0,32); mem_filters(6)(26) <= to_signed(0,32);
  mem_filters(6)(27) <= to_signed(0,32); mem_filters(6)(28) <= to_signed(0,32); mem_filters(6)(29) <= to_signed(0,32);
  mem_filters(6)(30) <= to_signed(0,32); mem_filters(6)(31) <= to_signed(0,32); mem_filters(6)(32) <= to_signed(0,32);
  mem_filters(6)(33) <= to_signed(0,32); mem_filters(6)(34) <= to_signed(0,32); mem_filters(6)(35) <= to_signed(0,32);
  mem_filters(6)(36) <= to_signed(0,32); mem_filters(6)(37) <= to_signed(0,32); mem_filters(6)(38) <= to_signed(0,32);
  mem_filters(6)(39) <= to_signed(0,32); mem_filters(6)(40) <= to_signed(0,32); mem_filters(6)(41) <= to_signed(0,32);
  mem_filters(6)(42) <= to_signed(0,32); mem_filters(6)(43) <= to_signed(0,32); mem_filters(6)(44) <= to_signed(0,32);
  mem_filters(6)(45) <= to_signed(0,32);
  mem_filters(6)(46) <= to_signed(0,32); mem_filters(6)(47) <= to_signed(0,32); mem_filters(6)(48) <= to_signed(0,32);
  mem_filters(6)(49) <= to_signed(0,32); mem_filters(6)(50) <= to_signed(0,32); mem_filters(6)(51) <= to_signed(0,32);
  mem_filters(6)(52) <= to_signed(0,32); mem_filters(6)(53) <= to_signed(0,32); mem_filters(6)(54) <= to_signed(0,32);
  mem_filters(6)(55) <= to_signed(0,32); mem_filters(6)(56) <= to_signed(0,32); mem_filters(6)(57) <= to_signed(0,32);
  mem_filters(6)(58) <= to_signed(0,32); mem_filters(6)(59) <= to_signed(0,32); mem_filters(6)(60) <= to_signed(0,32);
  mem_filters(6)(61) <= to_signed(0,32); mem_filters(6)(62) <= to_signed(0,32); mem_filters(6)(63) <= to_signed(0,32);
  mem_filters(6)(64) <= to_signed(0,32); mem_filters(6)(65) <= to_signed(0,32); mem_filters(6)(66) <= to_signed(0,32);
  mem_filters(6)(67) <= to_signed(0,32); mem_filters(6)(68) <= to_signed(0,32); mem_filters(6)(69) <= to_signed(0,32);
  mem_filters(6)(70) <= to_signed(0,32); mem_filters(6)(71) <= to_signed(0,32); mem_filters(6)(72) <= to_signed(0,32);
  mem_filters(6)(73) <= to_signed(0,32); mem_filters(6)(74) <= to_signed(0,32); mem_filters(6)(75) <= to_signed(0,32);
  mem_filters(6)(76) <= to_signed(0,32); mem_filters(6)(77) <= to_signed(0,32); mem_filters(6)(78) <= to_signed(0,32);
  mem_filters(6)(79) <= to_signed(0,32); mem_filters(6)(80) <= to_signed(0,32); mem_filters(6)(81) <= to_signed(0,32);
  mem_filters(6)(82) <= to_signed(0,32); mem_filters(6)(83) <= to_signed(0,32); mem_filters(6)(84) <= to_signed(0,32);
  mem_filters(6)(85) <= to_signed(0,32); mem_filters(6)(86) <= to_signed(0,32); mem_filters(6)(87) <= to_signed(0,32);
  mem_filters(6)(88) <= to_signed(0,32); mem_filters(6)(89) <= to_signed(0,32); mem_filters(6)(90) <= to_signed(0,32);
  mem_filters(6)(91) <= to_signed(0,32); mem_filters(6)(92) <= to_signed(0,32); mem_filters(6)(93) <= to_signed(0,32);
  mem_filters(6)(94) <= to_signed(0,32); mem_filters(6)(95) <= to_signed(0,32); mem_filters(6)(96) <= to_signed(0,32);
  mem_filters(6)(97) <= to_signed(0,32); mem_filters(6)(98) <= to_signed(0,32); mem_filters(6)(99) <= to_signed(0,32);
  mem_filters(6)(100) <= to_signed(0,32); mem_filters(6)(101) <= to_signed(0,32); mem_filters(6)(102) <= to_signed(0,32);
  mem_filters(6)(103) <= to_signed(0,32); mem_filters(6)(104) <= to_signed(0,32); mem_filters(6)(105) <= to_signed(0,32);
  mem_filters(6)(106) <= to_signed(0,32); mem_filters(6)(107) <= to_signed(0,32); mem_filters(6)(108) <= to_signed(0,32);
  mem_filters(6)(109) <= to_signed(0,32); mem_filters(6)(110) <= to_signed(0,32); mem_filters(6)(111) <= to_signed(0,32);
  mem_filters(6)(112) <= to_signed(0,32); mem_filters(6)(113) <= to_signed(0,32); mem_filters(6)(114) <= to_signed(0,32);
  mem_filters(6)(115) <= to_signed(0,32); mem_filters(6)(116) <= to_signed(0,32); mem_filters(6)(117) <= to_signed(0,32);
  mem_filters(6)(118) <= to_signed(0,32); mem_filters(6)(119) <= to_signed(0,32); mem_filters(6)(120) <= to_signed(0,32);
  mem_filters(6)(121) <= to_signed(0,32); mem_filters(6)(122) <= to_signed(0,32); mem_filters(6)(123) <= to_signed(0,32);
  mem_filters(6)(124) <= to_signed(0,32); mem_filters(6)(125) <= to_signed(0,32); mem_filters(6)(126) <= to_signed(0,32);
  mem_filters(6)(127) <= to_signed(0,32); mem_filters(6)(128) <= to_signed(0,32); mem_filters(6)(129) <= to_signed(0,32);
  mem_filters(6)(130) <= to_signed(0,32); mem_filters(6)(131) <= to_signed(0,32); mem_filters(6)(132) <= to_signed(0,32);
  mem_filters(6)(133) <= to_signed(0,32); mem_filters(6)(134) <= to_signed(0,32); mem_filters(6)(135) <= to_signed(0,32);
  mem_filters(6)(136) <= to_signed(0,32); mem_filters(6)(137) <= to_signed(0,32); mem_filters(6)(138) <= to_signed(0,32);
  mem_filters(6)(139) <= to_signed(0,32); mem_filters(6)(140) <= to_signed(0,32); mem_filters(6)(141) <= to_signed(0,32);
  mem_filters(6)(142) <= to_signed(0,32); mem_filters(6)(143) <= to_signed(0,32); mem_filters(6)(144) <= to_signed(0,32);
  mem_filters(6)(145) <= to_signed(0,32); mem_filters(6)(146) <= to_signed(0,32); mem_filters(6)(147) <= to_signed(0,32);
  mem_filters(6)(148) <= to_signed(0,32); mem_filters(6)(149) <= to_signed(0,32); mem_filters(6)(150) <= to_signed(0,32);
  mem_filters(6)(151) <= to_signed(0,32); mem_filters(6)(152) <= to_signed(0,32); mem_filters(6)(153) <= to_signed(0,32);
  mem_filters(6)(154) <= to_signed(0,32); mem_filters(6)(155) <= to_signed(0,32); mem_filters(6)(156) <= to_signed(0,32);
  mem_filters(6)(157) <= to_signed(0,32); mem_filters(6)(158) <= to_signed(0,32); mem_filters(6)(159) <= to_signed(0,32);
  mem_filters(6)(160) <= to_signed(0,32); mem_filters(6)(161) <= to_signed(0,32); mem_filters(6)(162) <= to_signed(0,32);
  mem_filters(6)(163) <= to_signed(0,32); mem_filters(6)(164) <= to_signed(0,32); mem_filters(6)(165) <= to_signed(0,32);
  mem_filters(6)(166) <= to_signed(0,32); mem_filters(6)(167) <= to_signed(0,32); mem_filters(6)(168) <= to_signed(0,32);
  mem_filters(6)(169) <= to_signed(0,32); mem_filters(6)(170) <= to_signed(0,32); mem_filters(6)(171) <= to_signed(0,32);
  mem_filters(6)(172) <= to_signed(0,32); mem_filters(6)(173) <= to_signed(0,32); mem_filters(6)(174) <= to_signed(0,32);
  mem_filters(6)(175) <= to_signed(0,32); mem_filters(6)(176) <= to_signed(0,32); mem_filters(6)(177) <= to_signed(0,32);
  mem_filters(6)(178) <= to_signed(0,32); mem_filters(6)(179) <= to_signed(0,32); mem_filters(6)(180) <= to_signed(0,32);
  mem_filters(6)(181) <= to_signed(0,32); mem_filters(6)(182) <= to_signed(0,32); mem_filters(6)(183) <= to_signed(0,32);
  mem_filters(6)(184) <= to_signed(0,32); mem_filters(6)(185) <= to_signed(0,32); mem_filters(6)(186) <= to_signed(0,32);
  mem_filters(6)(187) <= to_signed(0,32); mem_filters(6)(188) <= to_signed(0,32); mem_filters(6)(189) <= to_signed(0,32);
  mem_filters(6)(190) <= to_signed(0,32); mem_filters(6)(191) <= to_signed(0,32); mem_filters(6)(192) <= to_signed(0,32);
  mem_filters(6)(193) <= to_signed(0,32); mem_filters(6)(194) <= to_signed(0,32); mem_filters(6)(195) <= to_signed(0,32);
  mem_filters(6)(196) <= to_signed(0,32); mem_filters(6)(197) <= to_signed(0,32); mem_filters(6)(198) <= to_signed(0,32);
  mem_filters(6)(199) <= to_signed(0,32); mem_filters(6)(200) <= to_signed(0,32); mem_filters(6)(201) <= to_signed(0,32);
  mem_filters(6)(202) <= to_signed(0,32); mem_filters(6)(203) <= to_signed(0,32); mem_filters(6)(204) <= to_signed(0,32);
  mem_filters(6)(205) <= to_signed(0,32); mem_filters(6)(206) <= to_signed(0,32); mem_filters(6)(207) <= to_signed(0,32);
  mem_filters(6)(208) <= to_signed(0,32); mem_filters(6)(209) <= to_signed(0,32); mem_filters(6)(210) <= to_signed(0,32);
  mem_filters(6)(211) <= to_signed(0,32); mem_filters(6)(212) <= to_signed(0,32); mem_filters(6)(213) <= to_signed(0,32);
  mem_filters(6)(214) <= to_signed(0,32); mem_filters(6)(215) <= to_signed(0,32); mem_filters(6)(216) <= to_signed(0,32);
  mem_filters(6)(217) <= to_signed(0,32); mem_filters(6)(218) <= to_signed(0,32); mem_filters(6)(219) <= to_signed(0,32);
  mem_filters(6)(220) <= to_signed(0,32); mem_filters(6)(221) <= to_signed(0,32); mem_filters(6)(222) <= to_signed(0,32);
  mem_filters(6)(223) <= to_signed(0,32); mem_filters(6)(224) <= to_signed(0,32); mem_filters(6)(225) <= to_signed(0,32);
  mem_filters(6)(226) <= to_signed(0,32); mem_filters(6)(227) <= to_signed(0,32); mem_filters(6)(228) <= to_signed(0,32);
  mem_filters(6)(229) <= to_signed(0,32); mem_filters(6)(230) <= to_signed(0,32); mem_filters(6)(231) <= to_signed(0,32);
  mem_filters(6)(232) <= to_signed(0,32); mem_filters(6)(233) <= to_signed(0,32); mem_filters(6)(234) <= to_signed(0,32);
  mem_filters(6)(235) <= to_signed(0,32); mem_filters(6)(236) <= to_signed(0,32); mem_filters(6)(237) <= to_signed(0,32);
  mem_filters(6)(238) <= to_signed(0,32); mem_filters(6)(239) <= to_signed(0,32); mem_filters(6)(240) <= to_signed(0,32);
  mem_filters(6)(241) <= to_signed(0,32); mem_filters(6)(242) <= to_signed(0,32); mem_filters(6)(243) <= to_signed(0,32);
  mem_filters(6)(244) <= to_signed(0,32); mem_filters(6)(245) <= to_signed(0,32); mem_filters(6)(246) <= to_signed(0,32);
  mem_filters(6)(247) <= to_signed(0,32); mem_filters(6)(248) <= to_signed(0,32); mem_filters(6)(249) <= to_signed(0,32);
  mem_filters(6)(250) <= to_signed(0,32); mem_filters(6)(251) <= to_signed(0,32); mem_filters(6)(252) <= to_signed(0,32);
  mem_filters(6)(253) <= to_signed(0,32); mem_filters(6)(254) <= to_signed(0,32); mem_filters(6)(255) <= to_signed(0,32);
  
  --Filter 7
  mem_filters(7)(0) <= to_signed(0,32); mem_filters(7)(1) <= to_signed(0,32); mem_filters(7)(2) <= to_signed(0,32);
  mem_filters(7)(3) <= to_signed(0,32); mem_filters(7)(4) <= to_signed(0,32); mem_filters(7)(5) <= to_signed(0,32);
  mem_filters(7)(6) <= to_signed(0,32); mem_filters(7)(7) <= to_signed(0,32); mem_filters(7)(8) <= to_signed(0,32);
  mem_filters(7)(9) <= to_signed(0,32); mem_filters(7)(10) <= to_signed(0,32); mem_filters(7)(11) <= to_signed(0,32);
  mem_filters(7)(12) <= to_signed(0,32); mem_filters(7)(13) <= to_signed(0,32); mem_filters(7)(14) <= to_signed(0,32);
  mem_filters(7)(15) <= to_signed(0,32); mem_filters(7)(16) <= to_signed(0,32); mem_filters(7)(17) <= to_signed(0,32);
  mem_filters(7)(18) <= to_signed(0,32); mem_filters(7)(19) <= to_signed(0,32); mem_filters(7)(20) <= to_signed(0,32);
  mem_filters(7)(21) <= to_signed(0,32); mem_filters(7)(22) <= to_signed(0,32); mem_filters(7)(23) <= to_signed(0,32);
  mem_filters(7)(24) <= to_signed(0,32); mem_filters(7)(25) <= to_signed(0,32); mem_filters(7)(26) <= to_signed(0,32);
  mem_filters(7)(27) <= to_signed(0,32); mem_filters(7)(28) <= to_signed(0,32); mem_filters(7)(29) <= to_signed(0,32);
  mem_filters(7)(30) <= to_signed(0,32); mem_filters(7)(31) <= to_signed(0,32); mem_filters(7)(32) <= to_signed(0,32);
  mem_filters(7)(33) <= to_signed(0,32); mem_filters(7)(34) <= to_signed(0,32); mem_filters(7)(35) <= to_signed(0,32);
  mem_filters(7)(36) <= to_signed(0,32); mem_filters(7)(37) <= to_signed(0,32); mem_filters(7)(38) <= to_signed(0,32);
  mem_filters(7)(39) <= to_signed(0,32); mem_filters(7)(40) <= to_signed(0,32); mem_filters(7)(41) <= to_signed(0,32);
  mem_filters(7)(42) <= to_signed(0,32); mem_filters(7)(43) <= to_signed(0,32); mem_filters(7)(44) <= to_signed(0,32);
  mem_filters(7)(45) <= to_signed(0,32);
  mem_filters(7)(46) <= to_signed(0,32); mem_filters(7)(47) <= to_signed(0,32); mem_filters(7)(48) <= to_signed(0,32);
  mem_filters(7)(49) <= to_signed(0,32); mem_filters(7)(50) <= to_signed(0,32); mem_filters(7)(51) <= to_signed(0,32);
  mem_filters(7)(52) <= to_signed(0,32); mem_filters(7)(53) <= to_signed(0,32); mem_filters(7)(54) <= to_signed(0,32);
  mem_filters(7)(55) <= to_signed(0,32); mem_filters(7)(56) <= to_signed(0,32); mem_filters(7)(57) <= to_signed(0,32);
  mem_filters(7)(58) <= to_signed(0,32); mem_filters(7)(59) <= to_signed(0,32); mem_filters(7)(60) <= to_signed(0,32);
  mem_filters(7)(61) <= to_signed(0,32); mem_filters(7)(62) <= to_signed(0,32); mem_filters(7)(63) <= to_signed(0,32);
  mem_filters(7)(64) <= to_signed(0,32); mem_filters(7)(65) <= to_signed(0,32); mem_filters(7)(66) <= to_signed(0,32);
  mem_filters(7)(67) <= to_signed(0,32); mem_filters(7)(68) <= to_signed(0,32); mem_filters(7)(69) <= to_signed(0,32);
  mem_filters(7)(70) <= to_signed(0,32); mem_filters(7)(71) <= to_signed(0,32); mem_filters(7)(72) <= to_signed(0,32);
  mem_filters(7)(73) <= to_signed(0,32); mem_filters(7)(74) <= to_signed(0,32); mem_filters(7)(75) <= to_signed(0,32);
  mem_filters(7)(76) <= to_signed(0,32); mem_filters(7)(77) <= to_signed(0,32); mem_filters(7)(78) <= to_signed(0,32);
  mem_filters(7)(79) <= to_signed(0,32); mem_filters(7)(80) <= to_signed(0,32); mem_filters(7)(81) <= to_signed(0,32);
  mem_filters(7)(82) <= to_signed(0,32); mem_filters(7)(83) <= to_signed(0,32); mem_filters(7)(84) <= to_signed(0,32);
  mem_filters(7)(85) <= to_signed(0,32); mem_filters(7)(86) <= to_signed(0,32); mem_filters(7)(87) <= to_signed(0,32);
  mem_filters(7)(88) <= to_signed(0,32); mem_filters(7)(89) <= to_signed(0,32); mem_filters(7)(90) <= to_signed(0,32);
  mem_filters(7)(91) <= to_signed(0,32); mem_filters(7)(92) <= to_signed(0,32); mem_filters(7)(93) <= to_signed(0,32);
  mem_filters(7)(94) <= to_signed(0,32); mem_filters(7)(95) <= to_signed(0,32); mem_filters(7)(96) <= to_signed(0,32);
  mem_filters(7)(97) <= to_signed(0,32); mem_filters(7)(98) <= to_signed(0,32); mem_filters(7)(99) <= to_signed(0,32);
  mem_filters(7)(100) <= to_signed(0,32); mem_filters(7)(101) <= to_signed(0,32); mem_filters(7)(102) <= to_signed(0,32);
  mem_filters(7)(103) <= to_signed(0,32); mem_filters(7)(104) <= to_signed(0,32); mem_filters(7)(105) <= to_signed(0,32);
  mem_filters(7)(106) <= to_signed(0,32); mem_filters(7)(107) <= to_signed(0,32); mem_filters(7)(108) <= to_signed(0,32);
  mem_filters(7)(109) <= to_signed(0,32); mem_filters(7)(110) <= to_signed(0,32); mem_filters(7)(111) <= to_signed(0,32);
  mem_filters(7)(112) <= to_signed(0,32); mem_filters(7)(113) <= to_signed(0,32); mem_filters(7)(114) <= to_signed(0,32);
  mem_filters(7)(115) <= to_signed(0,32); mem_filters(7)(116) <= to_signed(0,32); mem_filters(7)(117) <= to_signed(0,32);
  mem_filters(7)(118) <= to_signed(0,32); mem_filters(7)(119) <= to_signed(0,32); mem_filters(7)(120) <= to_signed(0,32);
  mem_filters(7)(121) <= to_signed(0,32); mem_filters(7)(122) <= to_signed(0,32); mem_filters(7)(123) <= to_signed(0,32);
  mem_filters(7)(124) <= to_signed(0,32); mem_filters(7)(125) <= to_signed(0,32); mem_filters(7)(126) <= to_signed(0,32);
  mem_filters(7)(127) <= to_signed(0,32); mem_filters(7)(128) <= to_signed(0,32); mem_filters(7)(129) <= to_signed(0,32);
  mem_filters(7)(130) <= to_signed(0,32); mem_filters(7)(131) <= to_signed(0,32); mem_filters(7)(132) <= to_signed(0,32);
  mem_filters(7)(133) <= to_signed(0,32); mem_filters(7)(134) <= to_signed(0,32); mem_filters(7)(135) <= to_signed(0,32);
  mem_filters(7)(136) <= to_signed(0,32); mem_filters(7)(137) <= to_signed(0,32); mem_filters(7)(138) <= to_signed(0,32);
  mem_filters(7)(139) <= to_signed(0,32); mem_filters(7)(140) <= to_signed(0,32); mem_filters(7)(141) <= to_signed(0,32);
  mem_filters(7)(142) <= to_signed(0,32); mem_filters(7)(143) <= to_signed(0,32); mem_filters(7)(144) <= to_signed(0,32);
  mem_filters(7)(145) <= to_signed(0,32); mem_filters(7)(146) <= to_signed(0,32); mem_filters(7)(147) <= to_signed(0,32);
  mem_filters(7)(148) <= to_signed(0,32); mem_filters(7)(149) <= to_signed(0,32); mem_filters(7)(150) <= to_signed(0,32);
  mem_filters(7)(151) <= to_signed(0,32); mem_filters(7)(152) <= to_signed(0,32); mem_filters(7)(153) <= to_signed(0,32);
  mem_filters(7)(154) <= to_signed(0,32); mem_filters(7)(155) <= to_signed(0,32); mem_filters(7)(156) <= to_signed(0,32);
  mem_filters(7)(157) <= to_signed(0,32); mem_filters(7)(158) <= to_signed(0,32); mem_filters(7)(159) <= to_signed(0,32);
  mem_filters(7)(160) <= to_signed(0,32); mem_filters(7)(161) <= to_signed(0,32); mem_filters(7)(162) <= to_signed(0,32);
  mem_filters(7)(163) <= to_signed(0,32); mem_filters(7)(164) <= to_signed(0,32); mem_filters(7)(165) <= to_signed(0,32);
  mem_filters(7)(166) <= to_signed(0,32); mem_filters(7)(167) <= to_signed(0,32); mem_filters(7)(168) <= to_signed(0,32);
  mem_filters(7)(169) <= to_signed(0,32); mem_filters(7)(170) <= to_signed(0,32); mem_filters(7)(171) <= to_signed(0,32);
  mem_filters(7)(172) <= to_signed(0,32); mem_filters(7)(173) <= to_signed(0,32); mem_filters(7)(174) <= to_signed(0,32);
  mem_filters(7)(175) <= to_signed(0,32); mem_filters(7)(176) <= to_signed(0,32); mem_filters(7)(177) <= to_signed(0,32);
  mem_filters(7)(178) <= to_signed(0,32); mem_filters(7)(179) <= to_signed(0,32); mem_filters(7)(180) <= to_signed(0,32);
  mem_filters(7)(181) <= to_signed(0,32); mem_filters(7)(182) <= to_signed(0,32); mem_filters(7)(183) <= to_signed(0,32);
  mem_filters(7)(184) <= to_signed(0,32); mem_filters(7)(185) <= to_signed(0,32); mem_filters(7)(186) <= to_signed(0,32);
  mem_filters(7)(187) <= to_signed(0,32); mem_filters(7)(188) <= to_signed(0,32); mem_filters(7)(189) <= to_signed(0,32);
  mem_filters(7)(190) <= to_signed(0,32); mem_filters(7)(191) <= to_signed(0,32); mem_filters(7)(192) <= to_signed(0,32);
  mem_filters(7)(193) <= to_signed(0,32); mem_filters(7)(194) <= to_signed(0,32); mem_filters(7)(195) <= to_signed(0,32);
  mem_filters(7)(196) <= to_signed(0,32); mem_filters(7)(197) <= to_signed(0,32); mem_filters(7)(198) <= to_signed(0,32);
  mem_filters(7)(199) <= to_signed(0,32); mem_filters(7)(200) <= to_signed(0,32); mem_filters(7)(201) <= to_signed(0,32);
  mem_filters(7)(202) <= to_signed(0,32); mem_filters(7)(203) <= to_signed(0,32); mem_filters(7)(204) <= to_signed(0,32);
  mem_filters(7)(205) <= to_signed(0,32); mem_filters(7)(206) <= to_signed(0,32); mem_filters(7)(207) <= to_signed(0,32);
  mem_filters(7)(208) <= to_signed(0,32); mem_filters(7)(209) <= to_signed(0,32); mem_filters(7)(210) <= to_signed(0,32);
  mem_filters(7)(211) <= to_signed(0,32); mem_filters(7)(212) <= to_signed(0,32); mem_filters(7)(213) <= to_signed(0,32);
  mem_filters(7)(214) <= to_signed(0,32); mem_filters(7)(215) <= to_signed(0,32); mem_filters(7)(216) <= to_signed(0,32);
  mem_filters(7)(217) <= to_signed(0,32); mem_filters(7)(218) <= to_signed(0,32); mem_filters(7)(219) <= to_signed(0,32);
  mem_filters(7)(220) <= to_signed(0,32); mem_filters(7)(221) <= to_signed(0,32); mem_filters(7)(222) <= to_signed(0,32);
  mem_filters(7)(223) <= to_signed(0,32); mem_filters(7)(224) <= to_signed(0,32); mem_filters(7)(225) <= to_signed(0,32);
  mem_filters(7)(226) <= to_signed(0,32); mem_filters(7)(227) <= to_signed(0,32); mem_filters(7)(228) <= to_signed(0,32);
  mem_filters(7)(229) <= to_signed(0,32); mem_filters(7)(230) <= to_signed(0,32); mem_filters(7)(231) <= to_signed(0,32);
  mem_filters(7)(232) <= to_signed(0,32); mem_filters(7)(233) <= to_signed(0,32); mem_filters(7)(234) <= to_signed(0,32);
  mem_filters(7)(235) <= to_signed(0,32); mem_filters(7)(236) <= to_signed(0,32); mem_filters(7)(237) <= to_signed(0,32);
  mem_filters(7)(238) <= to_signed(0,32); mem_filters(7)(239) <= to_signed(0,32); mem_filters(7)(240) <= to_signed(0,32);
  mem_filters(7)(241) <= to_signed(0,32); mem_filters(7)(242) <= to_signed(0,32); mem_filters(7)(243) <= to_signed(0,32);
  mem_filters(7)(244) <= to_signed(0,32); mem_filters(7)(245) <= to_signed(0,32); mem_filters(7)(246) <= to_signed(0,32);
  mem_filters(7)(247) <= to_signed(0,32); mem_filters(7)(248) <= to_signed(0,32); mem_filters(7)(249) <= to_signed(0,32);
  mem_filters(7)(250) <= to_signed(0,32); mem_filters(7)(251) <= to_signed(0,32); mem_filters(7)(252) <= to_signed(0,32);
  mem_filters(7)(253) <= to_signed(0,32); mem_filters(7)(254) <= to_signed(0,32); mem_filters(7)(255) <= to_signed(0,32);
  
  --Filter 8
  mem_filters(8)(0) <= to_signed(0,32); mem_filters(8)(1) <= to_signed(0,32); mem_filters(8)(2) <= to_signed(0,32);
  mem_filters(8)(3) <= to_signed(0,32); mem_filters(8)(4) <= to_signed(0,32); mem_filters(8)(5) <= to_signed(0,32);
  mem_filters(8)(6) <= to_signed(0,32); mem_filters(8)(7) <= to_signed(0,32); mem_filters(8)(8) <= to_signed(0,32);
  mem_filters(8)(9) <= to_signed(0,32); mem_filters(8)(10) <= to_signed(0,32); mem_filters(8)(11) <= to_signed(0,32);
  mem_filters(8)(12) <= to_signed(0,32); mem_filters(8)(13) <= to_signed(0,32); mem_filters(8)(14) <= to_signed(0,32);
  mem_filters(8)(15) <= to_signed(0,32); mem_filters(8)(16) <= to_signed(0,32); mem_filters(8)(17) <= to_signed(0,32);
  mem_filters(8)(18) <= to_signed(0,32); mem_filters(8)(19) <= to_signed(0,32); mem_filters(8)(20) <= to_signed(0,32);
  mem_filters(8)(21) <= to_signed(0,32); mem_filters(8)(22) <= to_signed(0,32); mem_filters(8)(23) <= to_signed(0,32);
  mem_filters(8)(24) <= to_signed(0,32); mem_filters(8)(25) <= to_signed(0,32); mem_filters(8)(26) <= to_signed(0,32);
  mem_filters(8)(27) <= to_signed(0,32); mem_filters(8)(28) <= to_signed(0,32); mem_filters(8)(29) <= to_signed(0,32);
  mem_filters(8)(30) <= to_signed(0,32); mem_filters(8)(31) <= to_signed(0,32); mem_filters(8)(32) <= to_signed(0,32);
  mem_filters(8)(33) <= to_signed(0,32); mem_filters(8)(34) <= to_signed(0,32); mem_filters(8)(35) <= to_signed(0,32);
  mem_filters(8)(36) <= to_signed(0,32); mem_filters(8)(37) <= to_signed(0,32); mem_filters(8)(38) <= to_signed(0,32);
  mem_filters(8)(39) <= to_signed(0,32); mem_filters(8)(40) <= to_signed(0,32); mem_filters(8)(41) <= to_signed(0,32);
  mem_filters(8)(42) <= to_signed(0,32); mem_filters(8)(43) <= to_signed(0,32); mem_filters(8)(44) <= to_signed(0,32);
  mem_filters(8)(45) <= to_signed(0,32);
  mem_filters(8)(46) <= to_signed(0,32); mem_filters(8)(47) <= to_signed(0,32); mem_filters(8)(48) <= to_signed(0,32);
  mem_filters(8)(49) <= to_signed(0,32); mem_filters(8)(50) <= to_signed(0,32); mem_filters(8)(51) <= to_signed(0,32);
  mem_filters(8)(52) <= to_signed(0,32); mem_filters(8)(53) <= to_signed(0,32); mem_filters(8)(54) <= to_signed(0,32);
  mem_filters(8)(55) <= to_signed(0,32); mem_filters(8)(56) <= to_signed(0,32); mem_filters(8)(57) <= to_signed(0,32);
  mem_filters(8)(58) <= to_signed(0,32); mem_filters(8)(59) <= to_signed(0,32); mem_filters(8)(60) <= to_signed(0,32);
  mem_filters(8)(61) <= to_signed(0,32); mem_filters(8)(62) <= to_signed(0,32); mem_filters(8)(63) <= to_signed(0,32);
  mem_filters(8)(64) <= to_signed(0,32); mem_filters(8)(65) <= to_signed(0,32); mem_filters(8)(66) <= to_signed(0,32);
  mem_filters(8)(67) <= to_signed(0,32); mem_filters(8)(68) <= to_signed(0,32); mem_filters(8)(69) <= to_signed(0,32);
  mem_filters(8)(70) <= to_signed(0,32); mem_filters(8)(71) <= to_signed(0,32); mem_filters(8)(72) <= to_signed(0,32);
  mem_filters(8)(73) <= to_signed(0,32); mem_filters(8)(74) <= to_signed(0,32); mem_filters(8)(75) <= to_signed(0,32);
  mem_filters(8)(76) <= to_signed(0,32); mem_filters(8)(77) <= to_signed(0,32); mem_filters(8)(78) <= to_signed(0,32);
  mem_filters(8)(79) <= to_signed(0,32); mem_filters(8)(80) <= to_signed(0,32); mem_filters(8)(81) <= to_signed(0,32);
  mem_filters(8)(82) <= to_signed(0,32); mem_filters(8)(83) <= to_signed(0,32); mem_filters(8)(84) <= to_signed(0,32);
  mem_filters(8)(85) <= to_signed(0,32); mem_filters(8)(86) <= to_signed(0,32); mem_filters(8)(87) <= to_signed(0,32);
  mem_filters(8)(88) <= to_signed(0,32); mem_filters(8)(89) <= to_signed(0,32); mem_filters(8)(90) <= to_signed(0,32);
  mem_filters(8)(91) <= to_signed(0,32); mem_filters(8)(92) <= to_signed(0,32); mem_filters(8)(93) <= to_signed(0,32);
  mem_filters(8)(94) <= to_signed(0,32); mem_filters(8)(95) <= to_signed(0,32); mem_filters(8)(96) <= to_signed(0,32);
  mem_filters(8)(97) <= to_signed(0,32); mem_filters(8)(98) <= to_signed(0,32); mem_filters(8)(99) <= to_signed(0,32);
  mem_filters(8)(100) <= to_signed(0,32); mem_filters(8)(101) <= to_signed(0,32); mem_filters(8)(102) <= to_signed(0,32);
  mem_filters(8)(103) <= to_signed(0,32); mem_filters(8)(104) <= to_signed(0,32); mem_filters(8)(105) <= to_signed(0,32);
  mem_filters(8)(106) <= to_signed(0,32); mem_filters(8)(107) <= to_signed(0,32); mem_filters(8)(108) <= to_signed(0,32);
  mem_filters(8)(109) <= to_signed(0,32); mem_filters(8)(110) <= to_signed(0,32); mem_filters(8)(111) <= to_signed(0,32);
  mem_filters(8)(112) <= to_signed(0,32); mem_filters(8)(113) <= to_signed(0,32); mem_filters(8)(114) <= to_signed(0,32);
  mem_filters(8)(115) <= to_signed(0,32); mem_filters(8)(116) <= to_signed(0,32); mem_filters(8)(117) <= to_signed(0,32);
  mem_filters(8)(118) <= to_signed(0,32); mem_filters(8)(119) <= to_signed(0,32); mem_filters(8)(120) <= to_signed(0,32);
  mem_filters(8)(121) <= to_signed(0,32); mem_filters(8)(122) <= to_signed(0,32); mem_filters(8)(123) <= to_signed(0,32);
  mem_filters(8)(124) <= to_signed(0,32); mem_filters(8)(125) <= to_signed(0,32); mem_filters(8)(126) <= to_signed(0,32);
  mem_filters(8)(127) <= to_signed(0,32); mem_filters(8)(128) <= to_signed(0,32); mem_filters(8)(129) <= to_signed(0,32);
  mem_filters(8)(130) <= to_signed(0,32); mem_filters(8)(131) <= to_signed(0,32); mem_filters(8)(132) <= to_signed(0,32);
  mem_filters(8)(133) <= to_signed(0,32); mem_filters(8)(134) <= to_signed(0,32); mem_filters(8)(135) <= to_signed(0,32);
  mem_filters(8)(136) <= to_signed(0,32); mem_filters(8)(137) <= to_signed(0,32); mem_filters(8)(138) <= to_signed(0,32);
  mem_filters(8)(139) <= to_signed(0,32); mem_filters(8)(140) <= to_signed(0,32); mem_filters(8)(141) <= to_signed(0,32);
  mem_filters(8)(142) <= to_signed(0,32); mem_filters(8)(143) <= to_signed(0,32); mem_filters(8)(144) <= to_signed(0,32);
  mem_filters(8)(145) <= to_signed(0,32); mem_filters(8)(146) <= to_signed(0,32); mem_filters(8)(147) <= to_signed(0,32);
  mem_filters(8)(148) <= to_signed(0,32); mem_filters(8)(149) <= to_signed(0,32); mem_filters(8)(150) <= to_signed(0,32);
  mem_filters(8)(151) <= to_signed(0,32); mem_filters(8)(152) <= to_signed(0,32); mem_filters(8)(153) <= to_signed(0,32);
  mem_filters(8)(154) <= to_signed(0,32); mem_filters(8)(155) <= to_signed(0,32); mem_filters(8)(156) <= to_signed(0,32);
  mem_filters(8)(157) <= to_signed(0,32); mem_filters(8)(158) <= to_signed(0,32); mem_filters(8)(159) <= to_signed(0,32);
  mem_filters(8)(160) <= to_signed(0,32); mem_filters(8)(161) <= to_signed(0,32); mem_filters(8)(162) <= to_signed(0,32);
  mem_filters(8)(163) <= to_signed(0,32); mem_filters(8)(164) <= to_signed(0,32); mem_filters(8)(165) <= to_signed(0,32);
  mem_filters(8)(166) <= to_signed(0,32); mem_filters(8)(167) <= to_signed(0,32); mem_filters(8)(168) <= to_signed(0,32);
  mem_filters(8)(169) <= to_signed(0,32); mem_filters(8)(170) <= to_signed(0,32); mem_filters(8)(171) <= to_signed(0,32);
  mem_filters(8)(172) <= to_signed(0,32); mem_filters(8)(173) <= to_signed(0,32); mem_filters(8)(174) <= to_signed(0,32);
  mem_filters(8)(175) <= to_signed(0,32); mem_filters(8)(176) <= to_signed(0,32); mem_filters(8)(177) <= to_signed(0,32);
  mem_filters(8)(178) <= to_signed(0,32); mem_filters(8)(179) <= to_signed(0,32); mem_filters(8)(180) <= to_signed(0,32);
  mem_filters(8)(181) <= to_signed(0,32); mem_filters(8)(182) <= to_signed(0,32); mem_filters(8)(183) <= to_signed(0,32);
  mem_filters(8)(184) <= to_signed(0,32); mem_filters(8)(185) <= to_signed(0,32); mem_filters(8)(186) <= to_signed(0,32);
  mem_filters(8)(187) <= to_signed(0,32); mem_filters(8)(188) <= to_signed(0,32); mem_filters(8)(189) <= to_signed(0,32);
  mem_filters(8)(190) <= to_signed(0,32); mem_filters(8)(191) <= to_signed(0,32); mem_filters(8)(192) <= to_signed(0,32);
  mem_filters(8)(193) <= to_signed(0,32); mem_filters(8)(194) <= to_signed(0,32); mem_filters(8)(195) <= to_signed(0,32);
  mem_filters(8)(196) <= to_signed(0,32); mem_filters(8)(197) <= to_signed(0,32); mem_filters(8)(198) <= to_signed(0,32);
  mem_filters(8)(199) <= to_signed(0,32); mem_filters(8)(200) <= to_signed(0,32); mem_filters(8)(201) <= to_signed(0,32);
  mem_filters(8)(202) <= to_signed(0,32); mem_filters(8)(203) <= to_signed(0,32); mem_filters(8)(204) <= to_signed(0,32);
  mem_filters(8)(205) <= to_signed(0,32); mem_filters(8)(206) <= to_signed(0,32); mem_filters(8)(207) <= to_signed(0,32);
  mem_filters(8)(208) <= to_signed(0,32); mem_filters(8)(209) <= to_signed(0,32); mem_filters(8)(210) <= to_signed(0,32);
  mem_filters(8)(211) <= to_signed(0,32); mem_filters(8)(212) <= to_signed(0,32); mem_filters(8)(213) <= to_signed(0,32);
  mem_filters(8)(214) <= to_signed(0,32); mem_filters(8)(215) <= to_signed(0,32); mem_filters(8)(216) <= to_signed(0,32);
  mem_filters(8)(217) <= to_signed(0,32); mem_filters(8)(218) <= to_signed(0,32); mem_filters(8)(219) <= to_signed(0,32);
  mem_filters(8)(220) <= to_signed(0,32); mem_filters(8)(221) <= to_signed(0,32); mem_filters(8)(222) <= to_signed(0,32);
  mem_filters(8)(223) <= to_signed(0,32); mem_filters(8)(224) <= to_signed(0,32); mem_filters(8)(225) <= to_signed(0,32);
  mem_filters(8)(226) <= to_signed(0,32); mem_filters(8)(227) <= to_signed(0,32); mem_filters(8)(228) <= to_signed(0,32);
  mem_filters(8)(229) <= to_signed(0,32); mem_filters(8)(230) <= to_signed(0,32); mem_filters(8)(231) <= to_signed(0,32);
  mem_filters(8)(232) <= to_signed(0,32); mem_filters(8)(233) <= to_signed(0,32); mem_filters(8)(234) <= to_signed(0,32);
  mem_filters(8)(235) <= to_signed(0,32); mem_filters(8)(236) <= to_signed(0,32); mem_filters(8)(237) <= to_signed(0,32);
  mem_filters(8)(238) <= to_signed(0,32); mem_filters(8)(239) <= to_signed(0,32); mem_filters(8)(240) <= to_signed(0,32);
  mem_filters(8)(241) <= to_signed(0,32); mem_filters(8)(242) <= to_signed(0,32); mem_filters(8)(243) <= to_signed(0,32);
  mem_filters(8)(244) <= to_signed(0,32); mem_filters(8)(245) <= to_signed(0,32); mem_filters(8)(246) <= to_signed(0,32);
  mem_filters(8)(247) <= to_signed(0,32); mem_filters(8)(248) <= to_signed(0,32); mem_filters(8)(249) <= to_signed(0,32);
  mem_filters(8)(250) <= to_signed(0,32); mem_filters(8)(251) <= to_signed(0,32); mem_filters(8)(252) <= to_signed(0,32);
  mem_filters(8)(253) <= to_signed(0,32); mem_filters(8)(254) <= to_signed(0,32); mem_filters(8)(255) <= to_signed(0,32);
  
  --Filter 9
  mem_filters(9)(0) <= to_signed(0,32); mem_filters(9)(1) <= to_signed(0,32); mem_filters(9)(2) <= to_signed(0,32);
  mem_filters(9)(3) <= to_signed(0,32); mem_filters(9)(4) <= to_signed(0,32); mem_filters(9)(5) <= to_signed(0,32);
  mem_filters(9)(6) <= to_signed(0,32); mem_filters(9)(7) <= to_signed(0,32); mem_filters(9)(8) <= to_signed(0,32);
  mem_filters(9)(9) <= to_signed(0,32); mem_filters(9)(10) <= to_signed(0,32); mem_filters(9)(11) <= to_signed(0,32);
  mem_filters(9)(12) <= to_signed(0,32); mem_filters(9)(13) <= to_signed(0,32); mem_filters(9)(14) <= to_signed(0,32);
  mem_filters(9)(15) <= to_signed(0,32); mem_filters(9)(16) <= to_signed(0,32); mem_filters(9)(17) <= to_signed(0,32);
  mem_filters(9)(18) <= to_signed(0,32); mem_filters(9)(19) <= to_signed(0,32); mem_filters(9)(20) <= to_signed(0,32);
  mem_filters(9)(21) <= to_signed(0,32); mem_filters(9)(22) <= to_signed(0,32); mem_filters(9)(23) <= to_signed(0,32);
  mem_filters(9)(24) <= to_signed(0,32); mem_filters(9)(25) <= to_signed(0,32); mem_filters(9)(26) <= to_signed(0,32);
  mem_filters(9)(27) <= to_signed(0,32); mem_filters(9)(28) <= to_signed(0,32); mem_filters(9)(29) <= to_signed(0,32);
  mem_filters(9)(30) <= to_signed(0,32); mem_filters(9)(31) <= to_signed(0,32); mem_filters(9)(32) <= to_signed(0,32);
  mem_filters(9)(33) <= to_signed(0,32); mem_filters(9)(34) <= to_signed(0,32); mem_filters(9)(35) <= to_signed(0,32);
  mem_filters(9)(36) <= to_signed(0,32); mem_filters(9)(37) <= to_signed(0,32); mem_filters(9)(38) <= to_signed(0,32);
  mem_filters(9)(39) <= to_signed(0,32); mem_filters(9)(40) <= to_signed(0,32); mem_filters(9)(41) <= to_signed(0,32);
  mem_filters(9)(42) <= to_signed(0,32); mem_filters(9)(43) <= to_signed(0,32); mem_filters(9)(44) <= to_signed(0,32);
  mem_filters(9)(45) <= to_signed(0,32);
  mem_filters(9)(46) <= to_signed(0,32); mem_filters(9)(47) <= to_signed(0,32); mem_filters(9)(48) <= to_signed(0,32);
  mem_filters(9)(49) <= to_signed(0,32); mem_filters(9)(50) <= to_signed(0,32); mem_filters(9)(51) <= to_signed(0,32);
  mem_filters(9)(52) <= to_signed(0,32); mem_filters(9)(53) <= to_signed(0,32); mem_filters(9)(54) <= to_signed(0,32);
  mem_filters(9)(55) <= to_signed(0,32); mem_filters(9)(56) <= to_signed(0,32); mem_filters(9)(57) <= to_signed(0,32);
  mem_filters(9)(58) <= to_signed(0,32); mem_filters(9)(59) <= to_signed(0,32); mem_filters(9)(60) <= to_signed(0,32);
  mem_filters(9)(61) <= to_signed(0,32); mem_filters(9)(62) <= to_signed(0,32); mem_filters(9)(63) <= to_signed(0,32);
  mem_filters(9)(64) <= to_signed(0,32); mem_filters(9)(65) <= to_signed(0,32); mem_filters(9)(66) <= to_signed(0,32);
  mem_filters(9)(67) <= to_signed(0,32); mem_filters(9)(68) <= to_signed(0,32); mem_filters(9)(69) <= to_signed(0,32);
  mem_filters(9)(70) <= to_signed(0,32); mem_filters(9)(71) <= to_signed(0,32); mem_filters(9)(72) <= to_signed(0,32);
  mem_filters(9)(73) <= to_signed(0,32); mem_filters(9)(74) <= to_signed(0,32); mem_filters(9)(75) <= to_signed(0,32);
  mem_filters(9)(76) <= to_signed(0,32); mem_filters(9)(77) <= to_signed(0,32); mem_filters(9)(78) <= to_signed(0,32);
  mem_filters(9)(79) <= to_signed(0,32); mem_filters(9)(80) <= to_signed(0,32); mem_filters(9)(81) <= to_signed(0,32);
  mem_filters(9)(82) <= to_signed(0,32); mem_filters(9)(83) <= to_signed(0,32); mem_filters(9)(84) <= to_signed(0,32);
  mem_filters(9)(85) <= to_signed(0,32); mem_filters(9)(86) <= to_signed(0,32); mem_filters(9)(87) <= to_signed(0,32);
  mem_filters(9)(88) <= to_signed(0,32); mem_filters(9)(89) <= to_signed(0,32); mem_filters(9)(90) <= to_signed(0,32);
  mem_filters(9)(91) <= to_signed(0,32); mem_filters(9)(92) <= to_signed(0,32); mem_filters(9)(93) <= to_signed(0,32);
  mem_filters(9)(94) <= to_signed(0,32); mem_filters(9)(95) <= to_signed(0,32); mem_filters(9)(96) <= to_signed(0,32);
  mem_filters(9)(97) <= to_signed(0,32); mem_filters(9)(98) <= to_signed(0,32); mem_filters(9)(99) <= to_signed(0,32);
  mem_filters(9)(100) <= to_signed(0,32); mem_filters(9)(101) <= to_signed(0,32); mem_filters(9)(102) <= to_signed(0,32);
  mem_filters(9)(103) <= to_signed(0,32); mem_filters(9)(104) <= to_signed(0,32); mem_filters(9)(105) <= to_signed(0,32);
  mem_filters(9)(106) <= to_signed(0,32); mem_filters(9)(107) <= to_signed(0,32); mem_filters(9)(108) <= to_signed(0,32);
  mem_filters(9)(109) <= to_signed(0,32); mem_filters(9)(110) <= to_signed(0,32); mem_filters(9)(111) <= to_signed(0,32);
  mem_filters(9)(112) <= to_signed(0,32); mem_filters(9)(113) <= to_signed(0,32); mem_filters(9)(114) <= to_signed(0,32);
  mem_filters(9)(115) <= to_signed(0,32); mem_filters(9)(116) <= to_signed(0,32); mem_filters(9)(117) <= to_signed(0,32);
  mem_filters(9)(118) <= to_signed(0,32); mem_filters(9)(119) <= to_signed(0,32); mem_filters(9)(120) <= to_signed(0,32);
  mem_filters(9)(121) <= to_signed(0,32); mem_filters(9)(122) <= to_signed(0,32); mem_filters(9)(123) <= to_signed(0,32);
  mem_filters(9)(124) <= to_signed(0,32); mem_filters(9)(125) <= to_signed(0,32); mem_filters(9)(126) <= to_signed(0,32);
  mem_filters(9)(127) <= to_signed(0,32); mem_filters(9)(128) <= to_signed(0,32); mem_filters(9)(129) <= to_signed(0,32);
  mem_filters(9)(130) <= to_signed(0,32); mem_filters(9)(131) <= to_signed(0,32); mem_filters(9)(132) <= to_signed(0,32);
  mem_filters(9)(133) <= to_signed(0,32); mem_filters(9)(134) <= to_signed(0,32); mem_filters(9)(135) <= to_signed(0,32);
  mem_filters(9)(136) <= to_signed(0,32); mem_filters(9)(137) <= to_signed(0,32); mem_filters(9)(138) <= to_signed(0,32);
  mem_filters(9)(139) <= to_signed(0,32); mem_filters(9)(140) <= to_signed(0,32); mem_filters(9)(141) <= to_signed(0,32);
  mem_filters(9)(142) <= to_signed(0,32); mem_filters(9)(143) <= to_signed(0,32); mem_filters(9)(144) <= to_signed(0,32);
  mem_filters(9)(145) <= to_signed(0,32); mem_filters(9)(146) <= to_signed(0,32); mem_filters(9)(147) <= to_signed(0,32);
  mem_filters(9)(148) <= to_signed(0,32); mem_filters(9)(149) <= to_signed(0,32); mem_filters(9)(150) <= to_signed(0,32);
  mem_filters(9)(151) <= to_signed(0,32); mem_filters(9)(152) <= to_signed(0,32); mem_filters(9)(153) <= to_signed(0,32);
  mem_filters(9)(154) <= to_signed(0,32); mem_filters(9)(155) <= to_signed(0,32); mem_filters(9)(156) <= to_signed(0,32);
  mem_filters(9)(157) <= to_signed(0,32); mem_filters(9)(158) <= to_signed(0,32); mem_filters(9)(159) <= to_signed(0,32);
  mem_filters(9)(160) <= to_signed(0,32); mem_filters(9)(161) <= to_signed(0,32); mem_filters(9)(162) <= to_signed(0,32);
  mem_filters(9)(163) <= to_signed(0,32); mem_filters(9)(164) <= to_signed(0,32); mem_filters(9)(165) <= to_signed(0,32);
  mem_filters(9)(166) <= to_signed(0,32); mem_filters(9)(167) <= to_signed(0,32); mem_filters(9)(168) <= to_signed(0,32);
  mem_filters(9)(169) <= to_signed(0,32); mem_filters(9)(170) <= to_signed(0,32); mem_filters(9)(171) <= to_signed(0,32);
  mem_filters(9)(172) <= to_signed(0,32); mem_filters(9)(173) <= to_signed(0,32); mem_filters(9)(174) <= to_signed(0,32);
  mem_filters(9)(175) <= to_signed(0,32); mem_filters(9)(176) <= to_signed(0,32); mem_filters(9)(177) <= to_signed(0,32);
  mem_filters(9)(178) <= to_signed(0,32); mem_filters(9)(179) <= to_signed(0,32); mem_filters(9)(180) <= to_signed(0,32);
  mem_filters(9)(181) <= to_signed(0,32); mem_filters(9)(182) <= to_signed(0,32); mem_filters(9)(183) <= to_signed(0,32);
  mem_filters(9)(184) <= to_signed(0,32); mem_filters(9)(185) <= to_signed(0,32); mem_filters(9)(186) <= to_signed(0,32);
  mem_filters(9)(187) <= to_signed(0,32); mem_filters(9)(188) <= to_signed(0,32); mem_filters(9)(189) <= to_signed(0,32);
  mem_filters(9)(190) <= to_signed(0,32); mem_filters(9)(191) <= to_signed(0,32); mem_filters(9)(192) <= to_signed(0,32);
  mem_filters(9)(193) <= to_signed(0,32); mem_filters(9)(194) <= to_signed(0,32); mem_filters(9)(195) <= to_signed(0,32);
  mem_filters(9)(196) <= to_signed(0,32); mem_filters(9)(197) <= to_signed(0,32); mem_filters(9)(198) <= to_signed(0,32);
  mem_filters(9)(199) <= to_signed(0,32); mem_filters(9)(200) <= to_signed(0,32); mem_filters(9)(201) <= to_signed(0,32);
  mem_filters(9)(202) <= to_signed(0,32); mem_filters(9)(203) <= to_signed(0,32); mem_filters(9)(204) <= to_signed(0,32);
  mem_filters(9)(205) <= to_signed(0,32); mem_filters(9)(206) <= to_signed(0,32); mem_filters(9)(207) <= to_signed(0,32);
  mem_filters(9)(208) <= to_signed(0,32); mem_filters(9)(209) <= to_signed(0,32); mem_filters(9)(210) <= to_signed(0,32);
  mem_filters(9)(211) <= to_signed(0,32); mem_filters(9)(212) <= to_signed(0,32); mem_filters(9)(213) <= to_signed(0,32);
  mem_filters(9)(214) <= to_signed(0,32); mem_filters(9)(215) <= to_signed(0,32); mem_filters(9)(216) <= to_signed(0,32);
  mem_filters(9)(217) <= to_signed(0,32); mem_filters(9)(218) <= to_signed(0,32); mem_filters(9)(219) <= to_signed(0,32);
  mem_filters(9)(220) <= to_signed(0,32); mem_filters(9)(221) <= to_signed(0,32); mem_filters(9)(222) <= to_signed(0,32);
  mem_filters(9)(223) <= to_signed(0,32); mem_filters(9)(224) <= to_signed(0,32); mem_filters(9)(225) <= to_signed(0,32);
  mem_filters(9)(226) <= to_signed(0,32); mem_filters(9)(227) <= to_signed(0,32); mem_filters(9)(228) <= to_signed(0,32);
  mem_filters(9)(229) <= to_signed(0,32); mem_filters(9)(230) <= to_signed(0,32); mem_filters(9)(231) <= to_signed(0,32);
  mem_filters(9)(232) <= to_signed(0,32); mem_filters(9)(233) <= to_signed(0,32); mem_filters(9)(234) <= to_signed(0,32);
  mem_filters(9)(235) <= to_signed(0,32); mem_filters(9)(236) <= to_signed(0,32); mem_filters(9)(237) <= to_signed(0,32);
  mem_filters(9)(238) <= to_signed(0,32); mem_filters(9)(239) <= to_signed(0,32); mem_filters(9)(240) <= to_signed(0,32);
  mem_filters(9)(241) <= to_signed(0,32); mem_filters(9)(242) <= to_signed(0,32); mem_filters(9)(243) <= to_signed(0,32);
  mem_filters(9)(244) <= to_signed(0,32); mem_filters(9)(245) <= to_signed(0,32); mem_filters(9)(246) <= to_signed(0,32);
  mem_filters(9)(247) <= to_signed(0,32); mem_filters(9)(248) <= to_signed(0,32); mem_filters(9)(249) <= to_signed(0,32);
  mem_filters(9)(250) <= to_signed(0,32); mem_filters(9)(251) <= to_signed(0,32); mem_filters(9)(252) <= to_signed(0,32);
  mem_filters(9)(253) <= to_signed(0,32); mem_filters(9)(254) <= to_signed(0,32); mem_filters(9)(255) <= to_signed(0,32);
  
  --Filter 10
  mem_filters(10)(0) <= to_signed(0,32); mem_filters(10)(1) <= to_signed(0,32); mem_filters(10)(2) <= to_signed(0,32);
  mem_filters(10)(3) <= to_signed(0,32); mem_filters(10)(4) <= to_signed(0,32); mem_filters(10)(5) <= to_signed(0,32);
  mem_filters(10)(6) <= to_signed(0,32); mem_filters(10)(7) <= to_signed(0,32); mem_filters(10)(8) <= to_signed(0,32);
  mem_filters(10)(9) <= to_signed(0,32); mem_filters(10)(10) <= to_signed(0,32); mem_filters(10)(11) <= to_signed(0,32);
  mem_filters(10)(12) <= to_signed(0,32); mem_filters(10)(13) <= to_signed(0,32); mem_filters(10)(14) <= to_signed(0,32);
  mem_filters(10)(15) <= to_signed(0,32); mem_filters(10)(16) <= to_signed(0,32); mem_filters(10)(17) <= to_signed(0,32);
  mem_filters(10)(18) <= to_signed(0,32); mem_filters(10)(19) <= to_signed(0,32); mem_filters(10)(20) <= to_signed(0,32);
  mem_filters(10)(21) <= to_signed(0,32); mem_filters(10)(22) <= to_signed(0,32); mem_filters(10)(23) <= to_signed(0,32);
  mem_filters(10)(24) <= to_signed(0,32); mem_filters(10)(25) <= to_signed(0,32); mem_filters(10)(26) <= to_signed(0,32);
  mem_filters(10)(27) <= to_signed(0,32); mem_filters(10)(28) <= to_signed(0,32); mem_filters(10)(29) <= to_signed(0,32);
  mem_filters(10)(30) <= to_signed(0,32); mem_filters(10)(31) <= to_signed(0,32); mem_filters(10)(32) <= to_signed(0,32);
  mem_filters(10)(33) <= to_signed(0,32); mem_filters(10)(34) <= to_signed(0,32); mem_filters(10)(35) <= to_signed(0,32);
  mem_filters(10)(36) <= to_signed(0,32); mem_filters(10)(37) <= to_signed(0,32); mem_filters(10)(38) <= to_signed(0,32);
  mem_filters(10)(39) <= to_signed(0,32); mem_filters(10)(40) <= to_signed(0,32); mem_filters(10)(41) <= to_signed(0,32);
  mem_filters(10)(42) <= to_signed(0,32); mem_filters(10)(43) <= to_signed(0,32); mem_filters(10)(44) <= to_signed(0,32);
  mem_filters(10)(45) <= to_signed(0,32);
  mem_filters(10)(46) <= to_signed(0,32); mem_filters(10)(47) <= to_signed(0,32); mem_filters(10)(48) <= to_signed(0,32);
  mem_filters(10)(49) <= to_signed(0,32); mem_filters(10)(50) <= to_signed(0,32); mem_filters(10)(51) <= to_signed(0,32);
  mem_filters(10)(52) <= to_signed(0,32); mem_filters(10)(53) <= to_signed(0,32); mem_filters(10)(54) <= to_signed(0,32);
  mem_filters(10)(55) <= to_signed(0,32); mem_filters(10)(56) <= to_signed(0,32); mem_filters(10)(57) <= to_signed(0,32);
  mem_filters(10)(58) <= to_signed(0,32); mem_filters(10)(59) <= to_signed(0,32); mem_filters(10)(60) <= to_signed(0,32);
  mem_filters(10)(61) <= to_signed(0,32); mem_filters(10)(62) <= to_signed(0,32); mem_filters(10)(63) <= to_signed(0,32);
  mem_filters(10)(64) <= to_signed(0,32); mem_filters(10)(65) <= to_signed(0,32); mem_filters(10)(66) <= to_signed(0,32);
  mem_filters(10)(67) <= to_signed(0,32); mem_filters(10)(68) <= to_signed(0,32); mem_filters(10)(69) <= to_signed(0,32);
  mem_filters(10)(70) <= to_signed(0,32); mem_filters(10)(71) <= to_signed(0,32); mem_filters(10)(72) <= to_signed(0,32);
  mem_filters(10)(73) <= to_signed(0,32); mem_filters(10)(74) <= to_signed(0,32); mem_filters(10)(75) <= to_signed(0,32);
  mem_filters(10)(76) <= to_signed(0,32); mem_filters(10)(77) <= to_signed(0,32); mem_filters(10)(78) <= to_signed(0,32);
  mem_filters(10)(79) <= to_signed(0,32); mem_filters(10)(80) <= to_signed(0,32); mem_filters(10)(81) <= to_signed(0,32);
  mem_filters(10)(82) <= to_signed(0,32); mem_filters(10)(83) <= to_signed(0,32); mem_filters(10)(84) <= to_signed(0,32);
  mem_filters(10)(85) <= to_signed(0,32); mem_filters(10)(86) <= to_signed(0,32); mem_filters(10)(87) <= to_signed(0,32);
  mem_filters(10)(88) <= to_signed(0,32); mem_filters(10)(89) <= to_signed(0,32); mem_filters(10)(90) <= to_signed(0,32);
  mem_filters(10)(91) <= to_signed(0,32); mem_filters(10)(92) <= to_signed(0,32); mem_filters(10)(93) <= to_signed(0,32);
  mem_filters(10)(94) <= to_signed(0,32); mem_filters(10)(95) <= to_signed(0,32); mem_filters(10)(96) <= to_signed(0,32);
  mem_filters(10)(97) <= to_signed(0,32); mem_filters(10)(98) <= to_signed(0,32); mem_filters(10)(99) <= to_signed(0,32);
  mem_filters(10)(100) <= to_signed(0,32); mem_filters(10)(101) <= to_signed(0,32); mem_filters(10)(102) <= to_signed(0,32);
  mem_filters(10)(103) <= to_signed(0,32); mem_filters(10)(104) <= to_signed(0,32); mem_filters(10)(105) <= to_signed(0,32);
  mem_filters(10)(106) <= to_signed(0,32); mem_filters(10)(107) <= to_signed(0,32); mem_filters(10)(108) <= to_signed(0,32);
  mem_filters(10)(109) <= to_signed(0,32); mem_filters(10)(110) <= to_signed(0,32); mem_filters(10)(111) <= to_signed(0,32);
  mem_filters(10)(112) <= to_signed(0,32); mem_filters(10)(113) <= to_signed(0,32); mem_filters(10)(114) <= to_signed(0,32);
  mem_filters(10)(115) <= to_signed(0,32); mem_filters(10)(116) <= to_signed(0,32); mem_filters(10)(117) <= to_signed(0,32);
  mem_filters(10)(118) <= to_signed(0,32); mem_filters(10)(119) <= to_signed(0,32); mem_filters(10)(120) <= to_signed(0,32);
  mem_filters(10)(121) <= to_signed(0,32); mem_filters(10)(122) <= to_signed(0,32); mem_filters(10)(123) <= to_signed(0,32);
  mem_filters(10)(124) <= to_signed(0,32); mem_filters(10)(125) <= to_signed(0,32); mem_filters(10)(126) <= to_signed(0,32);
  mem_filters(10)(127) <= to_signed(0,32); mem_filters(10)(128) <= to_signed(0,32); mem_filters(10)(129) <= to_signed(0,32);
  mem_filters(10)(130) <= to_signed(0,32); mem_filters(10)(131) <= to_signed(0,32); mem_filters(10)(132) <= to_signed(0,32);
  mem_filters(10)(133) <= to_signed(0,32); mem_filters(10)(134) <= to_signed(0,32); mem_filters(10)(135) <= to_signed(0,32);
  mem_filters(10)(136) <= to_signed(0,32); mem_filters(10)(137) <= to_signed(0,32); mem_filters(10)(138) <= to_signed(0,32);
  mem_filters(10)(139) <= to_signed(0,32); mem_filters(10)(140) <= to_signed(0,32); mem_filters(10)(141) <= to_signed(0,32);
  mem_filters(10)(142) <= to_signed(0,32); mem_filters(10)(143) <= to_signed(0,32); mem_filters(10)(144) <= to_signed(0,32);
  mem_filters(10)(145) <= to_signed(0,32); mem_filters(10)(146) <= to_signed(0,32); mem_filters(10)(147) <= to_signed(0,32);
  mem_filters(10)(148) <= to_signed(0,32); mem_filters(10)(149) <= to_signed(0,32); mem_filters(10)(150) <= to_signed(0,32);
  mem_filters(10)(151) <= to_signed(0,32); mem_filters(10)(152) <= to_signed(0,32); mem_filters(10)(153) <= to_signed(0,32);
  mem_filters(10)(154) <= to_signed(0,32); mem_filters(10)(155) <= to_signed(0,32); mem_filters(10)(156) <= to_signed(0,32);
  mem_filters(10)(157) <= to_signed(0,32); mem_filters(10)(158) <= to_signed(0,32); mem_filters(10)(159) <= to_signed(0,32);
  mem_filters(10)(160) <= to_signed(0,32); mem_filters(10)(161) <= to_signed(0,32); mem_filters(10)(162) <= to_signed(0,32);
  mem_filters(10)(163) <= to_signed(0,32); mem_filters(10)(164) <= to_signed(0,32); mem_filters(10)(165) <= to_signed(0,32);
  mem_filters(10)(166) <= to_signed(0,32); mem_filters(10)(167) <= to_signed(0,32); mem_filters(10)(168) <= to_signed(0,32);
  mem_filters(10)(169) <= to_signed(0,32); mem_filters(10)(170) <= to_signed(0,32); mem_filters(10)(171) <= to_signed(0,32);
  mem_filters(10)(172) <= to_signed(0,32); mem_filters(10)(173) <= to_signed(0,32); mem_filters(10)(174) <= to_signed(0,32);
  mem_filters(10)(175) <= to_signed(0,32); mem_filters(10)(176) <= to_signed(0,32); mem_filters(10)(177) <= to_signed(0,32);
  mem_filters(10)(178) <= to_signed(0,32); mem_filters(10)(179) <= to_signed(0,32); mem_filters(10)(180) <= to_signed(0,32);
  mem_filters(10)(181) <= to_signed(0,32); mem_filters(10)(182) <= to_signed(0,32); mem_filters(10)(183) <= to_signed(0,32);
  mem_filters(10)(184) <= to_signed(0,32); mem_filters(10)(185) <= to_signed(0,32); mem_filters(10)(186) <= to_signed(0,32);
  mem_filters(10)(187) <= to_signed(0,32); mem_filters(10)(188) <= to_signed(0,32); mem_filters(10)(189) <= to_signed(0,32);
  mem_filters(10)(190) <= to_signed(0,32); mem_filters(10)(191) <= to_signed(0,32); mem_filters(10)(192) <= to_signed(0,32);
  mem_filters(10)(193) <= to_signed(0,32); mem_filters(10)(194) <= to_signed(0,32); mem_filters(10)(195) <= to_signed(0,32);
  mem_filters(10)(196) <= to_signed(0,32); mem_filters(10)(197) <= to_signed(0,32); mem_filters(10)(198) <= to_signed(0,32);
  mem_filters(10)(199) <= to_signed(0,32); mem_filters(10)(200) <= to_signed(0,32); mem_filters(10)(201) <= to_signed(0,32);
  mem_filters(10)(202) <= to_signed(0,32); mem_filters(10)(203) <= to_signed(0,32); mem_filters(10)(204) <= to_signed(0,32);
  mem_filters(10)(205) <= to_signed(0,32); mem_filters(10)(206) <= to_signed(0,32); mem_filters(10)(207) <= to_signed(0,32);
  mem_filters(10)(208) <= to_signed(0,32); mem_filters(10)(209) <= to_signed(0,32); mem_filters(10)(210) <= to_signed(0,32);
  mem_filters(10)(211) <= to_signed(0,32); mem_filters(10)(212) <= to_signed(0,32); mem_filters(10)(213) <= to_signed(0,32);
  mem_filters(10)(214) <= to_signed(0,32); mem_filters(10)(215) <= to_signed(0,32); mem_filters(10)(216) <= to_signed(0,32);
  mem_filters(10)(217) <= to_signed(0,32); mem_filters(10)(218) <= to_signed(0,32); mem_filters(10)(219) <= to_signed(0,32);
  mem_filters(10)(220) <= to_signed(0,32); mem_filters(10)(221) <= to_signed(0,32); mem_filters(10)(222) <= to_signed(0,32);
  mem_filters(10)(223) <= to_signed(0,32); mem_filters(10)(224) <= to_signed(0,32); mem_filters(10)(225) <= to_signed(0,32);
  mem_filters(10)(226) <= to_signed(0,32); mem_filters(10)(227) <= to_signed(0,32); mem_filters(10)(228) <= to_signed(0,32);
  mem_filters(10)(229) <= to_signed(0,32); mem_filters(10)(230) <= to_signed(0,32); mem_filters(10)(231) <= to_signed(0,32);
  mem_filters(10)(232) <= to_signed(0,32); mem_filters(10)(233) <= to_signed(0,32); mem_filters(10)(234) <= to_signed(0,32);
  mem_filters(10)(235) <= to_signed(0,32); mem_filters(10)(236) <= to_signed(0,32); mem_filters(10)(237) <= to_signed(0,32);
  mem_filters(10)(238) <= to_signed(0,32); mem_filters(10)(239) <= to_signed(0,32); mem_filters(10)(240) <= to_signed(0,32);
  mem_filters(10)(241) <= to_signed(0,32); mem_filters(10)(242) <= to_signed(0,32); mem_filters(10)(243) <= to_signed(0,32);
  mem_filters(10)(244) <= to_signed(0,32); mem_filters(10)(245) <= to_signed(0,32); mem_filters(10)(246) <= to_signed(0,32);
  mem_filters(10)(247) <= to_signed(0,32); mem_filters(10)(248) <= to_signed(0,32); mem_filters(10)(249) <= to_signed(0,32);
  mem_filters(10)(250) <= to_signed(0,32); mem_filters(10)(251) <= to_signed(0,32); mem_filters(10)(252) <= to_signed(0,32);
  mem_filters(10)(253) <= to_signed(0,32); mem_filters(10)(254) <= to_signed(0,32); mem_filters(10)(255) <= to_signed(0,32);
  
  --Filter 11
  mem_filters(11)(0) <= to_signed(0,32); mem_filters(11)(1) <= to_signed(0,32); mem_filters(11)(2) <= to_signed(0,32);
  mem_filters(11)(3) <= to_signed(0,32); mem_filters(11)(4) <= to_signed(0,32); mem_filters(11)(5) <= to_signed(0,32);
  mem_filters(11)(6) <= to_signed(0,32); mem_filters(11)(7) <= to_signed(0,32); mem_filters(11)(8) <= to_signed(0,32);
  mem_filters(11)(9) <= to_signed(0,32); mem_filters(11)(10) <= to_signed(0,32); mem_filters(11)(11) <= to_signed(0,32);
  mem_filters(11)(12) <= to_signed(0,32); mem_filters(11)(13) <= to_signed(0,32); mem_filters(11)(14) <= to_signed(0,32);
  mem_filters(11)(15) <= to_signed(0,32); mem_filters(11)(16) <= to_signed(0,32); mem_filters(11)(17) <= to_signed(0,32);
  mem_filters(11)(18) <= to_signed(0,32); mem_filters(11)(19) <= to_signed(0,32); mem_filters(11)(20) <= to_signed(0,32);
  mem_filters(11)(21) <= to_signed(0,32); mem_filters(11)(22) <= to_signed(0,32); mem_filters(11)(23) <= to_signed(0,32);
  mem_filters(11)(24) <= to_signed(0,32); mem_filters(11)(25) <= to_signed(0,32); mem_filters(11)(26) <= to_signed(0,32);
  mem_filters(11)(27) <= to_signed(0,32); mem_filters(11)(28) <= to_signed(0,32); mem_filters(11)(29) <= to_signed(0,32);
  mem_filters(11)(30) <= to_signed(0,32); mem_filters(11)(31) <= to_signed(0,32); mem_filters(11)(32) <= to_signed(0,32);
  mem_filters(11)(33) <= to_signed(0,32); mem_filters(11)(34) <= to_signed(0,32); mem_filters(11)(35) <= to_signed(0,32);
  mem_filters(11)(36) <= to_signed(0,32); mem_filters(11)(37) <= to_signed(0,32); mem_filters(11)(38) <= to_signed(0,32);
  mem_filters(11)(39) <= to_signed(0,32); mem_filters(11)(40) <= to_signed(0,32); mem_filters(11)(41) <= to_signed(0,32);
  mem_filters(11)(42) <= to_signed(0,32); mem_filters(11)(43) <= to_signed(0,32); mem_filters(11)(44) <= to_signed(0,32);
  mem_filters(11)(45) <= to_signed(0,32);
  mem_filters(11)(46) <= to_signed(0,32); mem_filters(11)(47) <= to_signed(0,32); mem_filters(11)(48) <= to_signed(0,32);
  mem_filters(11)(49) <= to_signed(0,32); mem_filters(11)(50) <= to_signed(0,32); mem_filters(11)(51) <= to_signed(0,32);
  mem_filters(11)(52) <= to_signed(0,32); mem_filters(11)(53) <= to_signed(0,32); mem_filters(11)(54) <= to_signed(0,32);
  mem_filters(11)(55) <= to_signed(0,32); mem_filters(11)(56) <= to_signed(0,32); mem_filters(11)(57) <= to_signed(0,32);
  mem_filters(11)(58) <= to_signed(0,32); mem_filters(11)(59) <= to_signed(0,32); mem_filters(11)(60) <= to_signed(0,32);
  mem_filters(11)(61) <= to_signed(0,32); mem_filters(11)(62) <= to_signed(0,32); mem_filters(11)(63) <= to_signed(0,32);
  mem_filters(11)(64) <= to_signed(0,32); mem_filters(11)(65) <= to_signed(0,32); mem_filters(11)(66) <= to_signed(0,32);
  mem_filters(11)(67) <= to_signed(0,32); mem_filters(11)(68) <= to_signed(0,32); mem_filters(11)(69) <= to_signed(0,32);
  mem_filters(11)(70) <= to_signed(0,32); mem_filters(11)(71) <= to_signed(0,32); mem_filters(11)(72) <= to_signed(0,32);
  mem_filters(11)(73) <= to_signed(0,32); mem_filters(11)(74) <= to_signed(0,32); mem_filters(11)(75) <= to_signed(0,32);
  mem_filters(11)(76) <= to_signed(0,32); mem_filters(11)(77) <= to_signed(0,32); mem_filters(11)(78) <= to_signed(0,32);
  mem_filters(11)(79) <= to_signed(0,32); mem_filters(11)(80) <= to_signed(0,32); mem_filters(11)(81) <= to_signed(0,32);
  mem_filters(11)(82) <= to_signed(0,32); mem_filters(11)(83) <= to_signed(0,32); mem_filters(11)(84) <= to_signed(0,32);
  mem_filters(11)(85) <= to_signed(0,32); mem_filters(11)(86) <= to_signed(0,32); mem_filters(11)(87) <= to_signed(0,32);
  mem_filters(11)(88) <= to_signed(0,32); mem_filters(11)(89) <= to_signed(0,32); mem_filters(11)(90) <= to_signed(0,32);
  mem_filters(11)(91) <= to_signed(0,32); mem_filters(11)(92) <= to_signed(0,32); mem_filters(11)(93) <= to_signed(0,32);
  mem_filters(11)(94) <= to_signed(0,32); mem_filters(11)(95) <= to_signed(0,32); mem_filters(11)(96) <= to_signed(0,32);
  mem_filters(11)(97) <= to_signed(0,32); mem_filters(11)(98) <= to_signed(0,32); mem_filters(11)(99) <= to_signed(0,32);
  mem_filters(11)(100) <= to_signed(0,32); mem_filters(11)(101) <= to_signed(0,32); mem_filters(11)(102) <= to_signed(0,32);
  mem_filters(11)(103) <= to_signed(0,32); mem_filters(11)(104) <= to_signed(0,32); mem_filters(11)(105) <= to_signed(0,32);
  mem_filters(11)(106) <= to_signed(0,32); mem_filters(11)(107) <= to_signed(0,32); mem_filters(11)(108) <= to_signed(0,32);
  mem_filters(11)(109) <= to_signed(0,32); mem_filters(11)(110) <= to_signed(0,32); mem_filters(11)(111) <= to_signed(0,32);
  mem_filters(11)(112) <= to_signed(0,32); mem_filters(11)(113) <= to_signed(0,32); mem_filters(11)(114) <= to_signed(0,32);
  mem_filters(11)(115) <= to_signed(0,32); mem_filters(11)(116) <= to_signed(0,32); mem_filters(11)(117) <= to_signed(0,32);
  mem_filters(11)(118) <= to_signed(0,32); mem_filters(11)(119) <= to_signed(0,32); mem_filters(11)(120) <= to_signed(0,32);
  mem_filters(11)(121) <= to_signed(0,32); mem_filters(11)(122) <= to_signed(0,32); mem_filters(11)(123) <= to_signed(0,32);
  mem_filters(11)(124) <= to_signed(0,32); mem_filters(11)(125) <= to_signed(0,32); mem_filters(11)(126) <= to_signed(0,32);
  mem_filters(11)(127) <= to_signed(0,32); mem_filters(11)(128) <= to_signed(0,32); mem_filters(11)(129) <= to_signed(0,32);
  mem_filters(11)(130) <= to_signed(0,32); mem_filters(11)(131) <= to_signed(0,32); mem_filters(11)(132) <= to_signed(0,32);
  mem_filters(11)(133) <= to_signed(0,32); mem_filters(11)(134) <= to_signed(0,32); mem_filters(11)(135) <= to_signed(0,32);
  mem_filters(11)(136) <= to_signed(0,32); mem_filters(11)(137) <= to_signed(0,32); mem_filters(11)(138) <= to_signed(0,32);
  mem_filters(11)(139) <= to_signed(0,32); mem_filters(11)(140) <= to_signed(0,32); mem_filters(11)(141) <= to_signed(0,32);
  mem_filters(11)(142) <= to_signed(0,32); mem_filters(11)(143) <= to_signed(0,32); mem_filters(11)(144) <= to_signed(0,32);
  mem_filters(11)(145) <= to_signed(0,32); mem_filters(11)(146) <= to_signed(0,32); mem_filters(11)(147) <= to_signed(0,32);
  mem_filters(11)(148) <= to_signed(0,32); mem_filters(11)(149) <= to_signed(0,32); mem_filters(11)(150) <= to_signed(0,32);
  mem_filters(11)(151) <= to_signed(0,32); mem_filters(11)(152) <= to_signed(0,32); mem_filters(11)(153) <= to_signed(0,32);
  mem_filters(11)(154) <= to_signed(0,32); mem_filters(11)(155) <= to_signed(0,32); mem_filters(11)(156) <= to_signed(0,32);
  mem_filters(11)(157) <= to_signed(0,32); mem_filters(11)(158) <= to_signed(0,32); mem_filters(11)(159) <= to_signed(0,32);
  mem_filters(11)(160) <= to_signed(0,32); mem_filters(11)(161) <= to_signed(0,32); mem_filters(11)(162) <= to_signed(0,32);
  mem_filters(11)(163) <= to_signed(0,32); mem_filters(11)(164) <= to_signed(0,32); mem_filters(11)(165) <= to_signed(0,32);
  mem_filters(11)(166) <= to_signed(0,32); mem_filters(11)(167) <= to_signed(0,32); mem_filters(11)(168) <= to_signed(0,32);
  mem_filters(11)(169) <= to_signed(0,32); mem_filters(11)(170) <= to_signed(0,32); mem_filters(11)(171) <= to_signed(0,32);
  mem_filters(11)(172) <= to_signed(0,32); mem_filters(11)(173) <= to_signed(0,32); mem_filters(11)(174) <= to_signed(0,32);
  mem_filters(11)(175) <= to_signed(0,32); mem_filters(11)(176) <= to_signed(0,32); mem_filters(11)(177) <= to_signed(0,32);
  mem_filters(11)(178) <= to_signed(0,32); mem_filters(11)(179) <= to_signed(0,32); mem_filters(11)(180) <= to_signed(0,32);
  mem_filters(11)(181) <= to_signed(0,32); mem_filters(11)(182) <= to_signed(0,32); mem_filters(11)(183) <= to_signed(0,32);
  mem_filters(11)(184) <= to_signed(0,32); mem_filters(11)(185) <= to_signed(0,32); mem_filters(11)(186) <= to_signed(0,32);
  mem_filters(11)(187) <= to_signed(0,32); mem_filters(11)(188) <= to_signed(0,32); mem_filters(11)(189) <= to_signed(0,32);
  mem_filters(11)(190) <= to_signed(0,32); mem_filters(11)(191) <= to_signed(0,32); mem_filters(11)(192) <= to_signed(0,32);
  mem_filters(11)(193) <= to_signed(0,32); mem_filters(11)(194) <= to_signed(0,32); mem_filters(11)(195) <= to_signed(0,32);
  mem_filters(11)(196) <= to_signed(0,32); mem_filters(11)(197) <= to_signed(0,32); mem_filters(11)(198) <= to_signed(0,32);
  mem_filters(11)(199) <= to_signed(0,32); mem_filters(11)(200) <= to_signed(0,32); mem_filters(11)(201) <= to_signed(0,32);
  mem_filters(11)(202) <= to_signed(0,32); mem_filters(11)(203) <= to_signed(0,32); mem_filters(11)(204) <= to_signed(0,32);
  mem_filters(11)(205) <= to_signed(0,32); mem_filters(11)(206) <= to_signed(0,32); mem_filters(11)(207) <= to_signed(0,32);
  mem_filters(11)(208) <= to_signed(0,32); mem_filters(11)(209) <= to_signed(0,32); mem_filters(11)(210) <= to_signed(0,32);
  mem_filters(11)(211) <= to_signed(0,32); mem_filters(11)(212) <= to_signed(0,32); mem_filters(11)(213) <= to_signed(0,32);
  mem_filters(11)(214) <= to_signed(0,32); mem_filters(11)(215) <= to_signed(0,32); mem_filters(11)(216) <= to_signed(0,32);
  mem_filters(11)(217) <= to_signed(0,32); mem_filters(11)(218) <= to_signed(0,32); mem_filters(11)(219) <= to_signed(0,32);
  mem_filters(11)(220) <= to_signed(0,32); mem_filters(11)(221) <= to_signed(0,32); mem_filters(11)(222) <= to_signed(0,32);
  mem_filters(11)(223) <= to_signed(0,32); mem_filters(11)(224) <= to_signed(0,32); mem_filters(11)(225) <= to_signed(0,32);
  mem_filters(11)(226) <= to_signed(0,32); mem_filters(11)(227) <= to_signed(0,32); mem_filters(11)(228) <= to_signed(0,32);
  mem_filters(11)(229) <= to_signed(0,32); mem_filters(11)(230) <= to_signed(0,32); mem_filters(11)(231) <= to_signed(0,32);
  mem_filters(11)(232) <= to_signed(0,32); mem_filters(11)(233) <= to_signed(0,32); mem_filters(11)(234) <= to_signed(0,32);
  mem_filters(11)(235) <= to_signed(0,32); mem_filters(11)(236) <= to_signed(0,32); mem_filters(11)(237) <= to_signed(0,32);
  mem_filters(11)(238) <= to_signed(0,32); mem_filters(11)(239) <= to_signed(0,32); mem_filters(11)(240) <= to_signed(0,32);
  mem_filters(11)(241) <= to_signed(0,32); mem_filters(11)(242) <= to_signed(0,32); mem_filters(11)(243) <= to_signed(0,32);
  mem_filters(11)(244) <= to_signed(0,32); mem_filters(11)(245) <= to_signed(0,32); mem_filters(11)(246) <= to_signed(0,32);
  mem_filters(11)(247) <= to_signed(0,32); mem_filters(11)(248) <= to_signed(0,32); mem_filters(11)(249) <= to_signed(0,32);
  mem_filters(11)(250) <= to_signed(0,32); mem_filters(11)(251) <= to_signed(0,32); mem_filters(11)(252) <= to_signed(0,32);
  mem_filters(11)(253) <= to_signed(0,32); mem_filters(11)(254) <= to_signed(0,32); mem_filters(11)(255) <= to_signed(0,32);
  
  --Filter 12
  mem_filters(12)(0) <= to_signed(0,32); mem_filters(12)(1) <= to_signed(0,32); mem_filters(12)(2) <= to_signed(0,32);
  mem_filters(12)(3) <= to_signed(0,32); mem_filters(12)(4) <= to_signed(0,32); mem_filters(12)(5) <= to_signed(0,32);
  mem_filters(12)(6) <= to_signed(0,32); mem_filters(12)(7) <= to_signed(0,32); mem_filters(12)(8) <= to_signed(0,32);
  mem_filters(12)(9) <= to_signed(0,32); mem_filters(12)(10) <= to_signed(0,32); mem_filters(12)(11) <= to_signed(0,32);
  mem_filters(12)(12) <= to_signed(0,32); mem_filters(12)(13) <= to_signed(0,32); mem_filters(12)(14) <= to_signed(0,32);
  mem_filters(12)(15) <= to_signed(0,32); mem_filters(12)(16) <= to_signed(0,32); mem_filters(12)(17) <= to_signed(0,32);
  mem_filters(12)(18) <= to_signed(0,32); mem_filters(12)(19) <= to_signed(0,32); mem_filters(12)(20) <= to_signed(0,32);
  mem_filters(12)(21) <= to_signed(0,32); mem_filters(12)(22) <= to_signed(0,32); mem_filters(12)(23) <= to_signed(0,32);
  mem_filters(12)(24) <= to_signed(0,32); mem_filters(12)(25) <= to_signed(0,32); mem_filters(12)(26) <= to_signed(0,32);
  mem_filters(12)(27) <= to_signed(0,32); mem_filters(12)(28) <= to_signed(0,32); mem_filters(12)(29) <= to_signed(0,32);
  mem_filters(12)(30) <= to_signed(0,32); mem_filters(12)(31) <= to_signed(0,32); mem_filters(12)(32) <= to_signed(0,32);
  mem_filters(12)(33) <= to_signed(0,32); mem_filters(12)(34) <= to_signed(0,32); mem_filters(12)(35) <= to_signed(0,32);
  mem_filters(12)(36) <= to_signed(0,32); mem_filters(12)(37) <= to_signed(0,32); mem_filters(12)(38) <= to_signed(0,32);
  mem_filters(12)(39) <= to_signed(0,32); mem_filters(12)(40) <= to_signed(0,32); mem_filters(12)(41) <= to_signed(0,32);
  mem_filters(12)(42) <= to_signed(0,32); mem_filters(12)(43) <= to_signed(0,32); mem_filters(12)(44) <= to_signed(0,32); 
  mem_filters(12)(45) <= to_signed(0,32);
  mem_filters(12)(46) <= to_signed(0,32); mem_filters(12)(47) <= to_signed(0,32); mem_filters(12)(48) <= to_signed(0,32);
  mem_filters(12)(49) <= to_signed(0,32); mem_filters(12)(50) <= to_signed(0,32); mem_filters(12)(51) <= to_signed(0,32);
  mem_filters(12)(52) <= to_signed(0,32); mem_filters(12)(53) <= to_signed(0,32); mem_filters(12)(54) <= to_signed(0,32);
  mem_filters(12)(55) <= to_signed(0,32); mem_filters(12)(56) <= to_signed(0,32); mem_filters(12)(57) <= to_signed(0,32);
  mem_filters(12)(58) <= to_signed(0,32); mem_filters(12)(59) <= to_signed(0,32); mem_filters(12)(60) <= to_signed(0,32);
  mem_filters(12)(61) <= to_signed(0,32); mem_filters(12)(62) <= to_signed(0,32); mem_filters(12)(63) <= to_signed(0,32);
  mem_filters(12)(64) <= to_signed(0,32); mem_filters(12)(65) <= to_signed(0,32); mem_filters(12)(66) <= to_signed(0,32);
  mem_filters(12)(67) <= to_signed(0,32); mem_filters(12)(68) <= to_signed(0,32); mem_filters(12)(69) <= to_signed(0,32);
  mem_filters(12)(70) <= to_signed(0,32); mem_filters(12)(71) <= to_signed(0,32); mem_filters(12)(72) <= to_signed(0,32);
  mem_filters(12)(73) <= to_signed(0,32); mem_filters(12)(74) <= to_signed(0,32); mem_filters(12)(75) <= to_signed(0,32);
  mem_filters(12)(76) <= to_signed(0,32); mem_filters(12)(77) <= to_signed(0,32); mem_filters(12)(78) <= to_signed(0,32);
  mem_filters(12)(79) <= to_signed(0,32); mem_filters(12)(80) <= to_signed(0,32); mem_filters(12)(81) <= to_signed(0,32);
  mem_filters(12)(82) <= to_signed(0,32); mem_filters(12)(83) <= to_signed(0,32); mem_filters(12)(84) <= to_signed(0,32);
  mem_filters(12)(85) <= to_signed(0,32); mem_filters(12)(86) <= to_signed(0,32); mem_filters(12)(87) <= to_signed(0,32);
  mem_filters(12)(88) <= to_signed(0,32); mem_filters(12)(89) <= to_signed(0,32); mem_filters(12)(90) <= to_signed(0,32);
  mem_filters(12)(91) <= to_signed(0,32); mem_filters(12)(92) <= to_signed(0,32); mem_filters(12)(93) <= to_signed(0,32);
  mem_filters(12)(94) <= to_signed(0,32); mem_filters(12)(95) <= to_signed(0,32); mem_filters(12)(96) <= to_signed(0,32);
  mem_filters(12)(97) <= to_signed(0,32); mem_filters(12)(98) <= to_signed(0,32); mem_filters(12)(99) <= to_signed(0,32);
  mem_filters(12)(100) <= to_signed(0,32); mem_filters(12)(101) <= to_signed(0,32); mem_filters(12)(102) <= to_signed(0,32);
  mem_filters(12)(103) <= to_signed(0,32); mem_filters(12)(104) <= to_signed(0,32); mem_filters(12)(105) <= to_signed(0,32);
  mem_filters(12)(106) <= to_signed(0,32); mem_filters(12)(107) <= to_signed(0,32); mem_filters(12)(108) <= to_signed(0,32);
  mem_filters(12)(109) <= to_signed(0,32); mem_filters(12)(110) <= to_signed(0,32); mem_filters(12)(111) <= to_signed(0,32);
  mem_filters(12)(112) <= to_signed(0,32); mem_filters(12)(113) <= to_signed(0,32); mem_filters(12)(114) <= to_signed(0,32);
  mem_filters(12)(115) <= to_signed(0,32); mem_filters(12)(116) <= to_signed(0,32); mem_filters(12)(117) <= to_signed(0,32);
  mem_filters(12)(118) <= to_signed(0,32); mem_filters(12)(119) <= to_signed(0,32); mem_filters(12)(120) <= to_signed(0,32);
  mem_filters(12)(121) <= to_signed(0,32); mem_filters(12)(122) <= to_signed(0,32); mem_filters(12)(123) <= to_signed(0,32);
  mem_filters(12)(124) <= to_signed(0,32); mem_filters(12)(125) <= to_signed(0,32); mem_filters(12)(126) <= to_signed(0,32);
  mem_filters(12)(127) <= to_signed(0,32); mem_filters(12)(128) <= to_signed(0,32); mem_filters(12)(129) <= to_signed(0,32);
  mem_filters(12)(130) <= to_signed(0,32); mem_filters(12)(131) <= to_signed(0,32); mem_filters(12)(132) <= to_signed(0,32);
  mem_filters(12)(133) <= to_signed(0,32); mem_filters(12)(134) <= to_signed(0,32); mem_filters(12)(135) <= to_signed(0,32);
  mem_filters(12)(136) <= to_signed(0,32); mem_filters(12)(137) <= to_signed(0,32); mem_filters(12)(138) <= to_signed(0,32);
  mem_filters(12)(139) <= to_signed(0,32); mem_filters(12)(140) <= to_signed(0,32); mem_filters(12)(141) <= to_signed(0,32);
  mem_filters(12)(142) <= to_signed(0,32); mem_filters(12)(143) <= to_signed(0,32); mem_filters(12)(144) <= to_signed(0,32);
  mem_filters(12)(145) <= to_signed(0,32); mem_filters(12)(146) <= to_signed(0,32); mem_filters(12)(147) <= to_signed(0,32);
  mem_filters(12)(148) <= to_signed(0,32); mem_filters(12)(149) <= to_signed(0,32); mem_filters(12)(150) <= to_signed(0,32);
  mem_filters(12)(151) <= to_signed(0,32); mem_filters(12)(152) <= to_signed(0,32); mem_filters(12)(153) <= to_signed(0,32);
  mem_filters(12)(154) <= to_signed(0,32); mem_filters(12)(155) <= to_signed(0,32); mem_filters(12)(156) <= to_signed(0,32);
  mem_filters(12)(157) <= to_signed(0,32); mem_filters(12)(158) <= to_signed(0,32); mem_filters(12)(159) <= to_signed(0,32);
  mem_filters(12)(160) <= to_signed(0,32); mem_filters(12)(161) <= to_signed(0,32); mem_filters(12)(162) <= to_signed(0,32);
  mem_filters(12)(163) <= to_signed(0,32); mem_filters(12)(164) <= to_signed(0,32); mem_filters(12)(165) <= to_signed(0,32);
  mem_filters(12)(166) <= to_signed(0,32); mem_filters(12)(167) <= to_signed(0,32); mem_filters(12)(168) <= to_signed(0,32);
  mem_filters(12)(169) <= to_signed(0,32); mem_filters(12)(170) <= to_signed(0,32); mem_filters(12)(171) <= to_signed(0,32);
  mem_filters(12)(172) <= to_signed(0,32); mem_filters(12)(173) <= to_signed(0,32); mem_filters(12)(174) <= to_signed(0,32);
  mem_filters(12)(175) <= to_signed(0,32); mem_filters(12)(176) <= to_signed(0,32); mem_filters(12)(177) <= to_signed(0,32);
  mem_filters(12)(178) <= to_signed(0,32); mem_filters(12)(179) <= to_signed(0,32); mem_filters(12)(180) <= to_signed(0,32);
  mem_filters(12)(181) <= to_signed(0,32); mem_filters(12)(182) <= to_signed(0,32); mem_filters(12)(183) <= to_signed(0,32);
  mem_filters(12)(184) <= to_signed(0,32); mem_filters(12)(185) <= to_signed(0,32); mem_filters(12)(186) <= to_signed(0,32);
  mem_filters(12)(187) <= to_signed(0,32); mem_filters(12)(188) <= to_signed(0,32); mem_filters(12)(189) <= to_signed(0,32);
  mem_filters(12)(190) <= to_signed(0,32); mem_filters(12)(191) <= to_signed(0,32); mem_filters(12)(192) <= to_signed(0,32);
  mem_filters(12)(193) <= to_signed(0,32); mem_filters(12)(194) <= to_signed(0,32); mem_filters(12)(195) <= to_signed(0,32);
  mem_filters(12)(196) <= to_signed(0,32); mem_filters(12)(197) <= to_signed(0,32); mem_filters(12)(198) <= to_signed(0,32);
  mem_filters(12)(199) <= to_signed(0,32); mem_filters(12)(200) <= to_signed(0,32); mem_filters(12)(201) <= to_signed(0,32);
  mem_filters(12)(202) <= to_signed(0,32); mem_filters(12)(203) <= to_signed(0,32); mem_filters(12)(204) <= to_signed(0,32);
  mem_filters(12)(205) <= to_signed(0,32); mem_filters(12)(206) <= to_signed(0,32); mem_filters(12)(207) <= to_signed(0,32);
  mem_filters(12)(208) <= to_signed(0,32); mem_filters(12)(209) <= to_signed(0,32); mem_filters(12)(210) <= to_signed(0,32);
  mem_filters(12)(211) <= to_signed(0,32); mem_filters(12)(212) <= to_signed(0,32); mem_filters(12)(213) <= to_signed(0,32);
  mem_filters(12)(214) <= to_signed(0,32); mem_filters(12)(215) <= to_signed(0,32); mem_filters(12)(216) <= to_signed(0,32);
  mem_filters(12)(217) <= to_signed(0,32); mem_filters(12)(218) <= to_signed(0,32); mem_filters(12)(219) <= to_signed(0,32);
  mem_filters(12)(220) <= to_signed(0,32); mem_filters(12)(221) <= to_signed(0,32); mem_filters(12)(222) <= to_signed(0,32);
  mem_filters(12)(223) <= to_signed(0,32); mem_filters(12)(224) <= to_signed(0,32); mem_filters(12)(225) <= to_signed(0,32);
  mem_filters(12)(226) <= to_signed(0,32); mem_filters(12)(227) <= to_signed(0,32); mem_filters(12)(228) <= to_signed(0,32);
  mem_filters(12)(229) <= to_signed(0,32); mem_filters(12)(230) <= to_signed(0,32); mem_filters(12)(231) <= to_signed(0,32);
  mem_filters(12)(232) <= to_signed(0,32); mem_filters(12)(233) <= to_signed(0,32); mem_filters(12)(234) <= to_signed(0,32);
  mem_filters(12)(235) <= to_signed(0,32); mem_filters(12)(236) <= to_signed(0,32); mem_filters(12)(237) <= to_signed(0,32);
  mem_filters(12)(238) <= to_signed(0,32); mem_filters(12)(239) <= to_signed(0,32); mem_filters(12)(240) <= to_signed(0,32);
  mem_filters(12)(241) <= to_signed(0,32); mem_filters(12)(242) <= to_signed(0,32); mem_filters(12)(243) <= to_signed(0,32);
  mem_filters(12)(244) <= to_signed(0,32); mem_filters(12)(245) <= to_signed(0,32); mem_filters(12)(246) <= to_signed(0,32);
  mem_filters(12)(247) <= to_signed(0,32); mem_filters(12)(248) <= to_signed(0,32); mem_filters(12)(249) <= to_signed(0,32);
  mem_filters(12)(250) <= to_signed(0,32); mem_filters(12)(251) <= to_signed(0,32); mem_filters(12)(252) <= to_signed(0,32);
  mem_filters(12)(253) <= to_signed(0,32); mem_filters(12)(254) <= to_signed(0,32); mem_filters(12)(255) <= to_signed(0,32);
  
  --Filter 13
  mem_filters(13)(0) <= to_signed(0,32); mem_filters(13)(1) <= to_signed(0,32); mem_filters(13)(2) <= to_signed(0,32);
  mem_filters(13)(3) <= to_signed(0,32); mem_filters(13)(4) <= to_signed(0,32); mem_filters(13)(5) <= to_signed(0,32);
  mem_filters(13)(6) <= to_signed(0,32); mem_filters(13)(7) <= to_signed(0,32); mem_filters(13)(8) <= to_signed(0,32);
  mem_filters(13)(9) <= to_signed(0,32); mem_filters(13)(10) <= to_signed(0,32); mem_filters(13)(11) <= to_signed(0,32);
  mem_filters(13)(12) <= to_signed(0,32); mem_filters(13)(13) <= to_signed(0,32); mem_filters(13)(14) <= to_signed(0,32);
  mem_filters(13)(15) <= to_signed(0,32); mem_filters(13)(16) <= to_signed(0,32); mem_filters(13)(17) <= to_signed(0,32);
  mem_filters(13)(18) <= to_signed(0,32); mem_filters(13)(19) <= to_signed(0,32); mem_filters(13)(20) <= to_signed(0,32);
  mem_filters(13)(21) <= to_signed(0,32); mem_filters(13)(22) <= to_signed(0,32); mem_filters(13)(23) <= to_signed(0,32);
  mem_filters(13)(24) <= to_signed(0,32); mem_filters(13)(25) <= to_signed(0,32); mem_filters(13)(26) <= to_signed(0,32);
  mem_filters(13)(27) <= to_signed(0,32); mem_filters(13)(28) <= to_signed(0,32); mem_filters(13)(29) <= to_signed(0,32);
  mem_filters(13)(30) <= to_signed(0,32); mem_filters(13)(31) <= to_signed(0,32); mem_filters(13)(32) <= to_signed(0,32);
  mem_filters(13)(33) <= to_signed(0,32); mem_filters(13)(34) <= to_signed(0,32); mem_filters(13)(35) <= to_signed(0,32);
  mem_filters(13)(36) <= to_signed(0,32); mem_filters(13)(37) <= to_signed(0,32); mem_filters(13)(38) <= to_signed(0,32);
  mem_filters(13)(39) <= to_signed(0,32); mem_filters(13)(40) <= to_signed(0,32); mem_filters(13)(41) <= to_signed(0,32);
  mem_filters(13)(42) <= to_signed(0,32); mem_filters(13)(43) <= to_signed(0,32); mem_filters(13)(44) <= to_signed(0,32);
  mem_filters(13)(45) <= to_signed(0,32);
  mem_filters(13)(46) <= to_signed(0,32); mem_filters(13)(47) <= to_signed(0,32); mem_filters(13)(48) <= to_signed(0,32);
  mem_filters(13)(49) <= to_signed(0,32); mem_filters(13)(50) <= to_signed(0,32); mem_filters(13)(51) <= to_signed(0,32);
  mem_filters(13)(52) <= to_signed(0,32); mem_filters(13)(53) <= to_signed(0,32); mem_filters(13)(54) <= to_signed(0,32);
  mem_filters(13)(55) <= to_signed(0,32); mem_filters(13)(56) <= to_signed(0,32); mem_filters(13)(57) <= to_signed(0,32);
  mem_filters(13)(58) <= to_signed(0,32); mem_filters(13)(59) <= to_signed(0,32); mem_filters(13)(60) <= to_signed(0,32);
  mem_filters(13)(61) <= to_signed(0,32); mem_filters(13)(62) <= to_signed(0,32); mem_filters(13)(63) <= to_signed(0,32);
  mem_filters(13)(64) <= to_signed(0,32); mem_filters(13)(65) <= to_signed(0,32); mem_filters(13)(66) <= to_signed(0,32);
  mem_filters(13)(67) <= to_signed(0,32); mem_filters(13)(68) <= to_signed(0,32); mem_filters(13)(69) <= to_signed(0,32);
  mem_filters(13)(70) <= to_signed(0,32); mem_filters(13)(71) <= to_signed(0,32); mem_filters(13)(72) <= to_signed(0,32);
  mem_filters(13)(73) <= to_signed(0,32); mem_filters(13)(74) <= to_signed(0,32); mem_filters(13)(75) <= to_signed(0,32);
  mem_filters(13)(76) <= to_signed(0,32); mem_filters(13)(77) <= to_signed(0,32); mem_filters(13)(78) <= to_signed(0,32);
  mem_filters(13)(79) <= to_signed(0,32); mem_filters(13)(80) <= to_signed(0,32); mem_filters(13)(81) <= to_signed(0,32);
  mem_filters(13)(82) <= to_signed(0,32); mem_filters(13)(83) <= to_signed(0,32); mem_filters(13)(84) <= to_signed(0,32);
  mem_filters(13)(85) <= to_signed(0,32); mem_filters(13)(86) <= to_signed(0,32); mem_filters(13)(87) <= to_signed(0,32);
  mem_filters(13)(88) <= to_signed(0,32); mem_filters(13)(89) <= to_signed(0,32); mem_filters(13)(90) <= to_signed(0,32);
  mem_filters(13)(91) <= to_signed(0,32); mem_filters(13)(92) <= to_signed(0,32); mem_filters(13)(93) <= to_signed(0,32);
  mem_filters(13)(94) <= to_signed(0,32); mem_filters(13)(95) <= to_signed(0,32); mem_filters(13)(96) <= to_signed(0,32);
  mem_filters(13)(97) <= to_signed(0,32); mem_filters(13)(98) <= to_signed(0,32); mem_filters(13)(99) <= to_signed(0,32);
  mem_filters(13)(100) <= to_signed(0,32); mem_filters(13)(101) <= to_signed(0,32); mem_filters(13)(102) <= to_signed(0,32);
  mem_filters(13)(103) <= to_signed(0,32); mem_filters(13)(104) <= to_signed(0,32); mem_filters(13)(105) <= to_signed(0,32);
  mem_filters(13)(106) <= to_signed(0,32); mem_filters(13)(107) <= to_signed(0,32); mem_filters(13)(108) <= to_signed(0,32);
  mem_filters(13)(109) <= to_signed(0,32); mem_filters(13)(110) <= to_signed(0,32); mem_filters(13)(111) <= to_signed(0,32);
  mem_filters(13)(112) <= to_signed(0,32); mem_filters(13)(113) <= to_signed(0,32); mem_filters(13)(114) <= to_signed(0,32);
  mem_filters(13)(115) <= to_signed(0,32); mem_filters(13)(116) <= to_signed(0,32); mem_filters(13)(117) <= to_signed(0,32);
  mem_filters(13)(118) <= to_signed(0,32); mem_filters(13)(119) <= to_signed(0,32); mem_filters(13)(120) <= to_signed(0,32);
  mem_filters(13)(121) <= to_signed(0,32); mem_filters(13)(122) <= to_signed(0,32); mem_filters(13)(123) <= to_signed(0,32);
  mem_filters(13)(124) <= to_signed(0,32); mem_filters(13)(125) <= to_signed(0,32); mem_filters(13)(126) <= to_signed(0,32);
  mem_filters(13)(127) <= to_signed(0,32); mem_filters(13)(128) <= to_signed(0,32); mem_filters(13)(129) <= to_signed(0,32);
  mem_filters(13)(130) <= to_signed(0,32); mem_filters(13)(131) <= to_signed(0,32); mem_filters(13)(132) <= to_signed(0,32);
  mem_filters(13)(133) <= to_signed(0,32); mem_filters(13)(134) <= to_signed(0,32); mem_filters(13)(135) <= to_signed(0,32);
  mem_filters(13)(136) <= to_signed(0,32); mem_filters(13)(137) <= to_signed(0,32); mem_filters(13)(138) <= to_signed(0,32);
  mem_filters(13)(139) <= to_signed(0,32); mem_filters(13)(140) <= to_signed(0,32); mem_filters(13)(141) <= to_signed(0,32);
  mem_filters(13)(142) <= to_signed(0,32); mem_filters(13)(143) <= to_signed(0,32); mem_filters(13)(144) <= to_signed(0,32);
  mem_filters(13)(145) <= to_signed(0,32); mem_filters(13)(146) <= to_signed(0,32); mem_filters(13)(147) <= to_signed(0,32);
  mem_filters(13)(148) <= to_signed(0,32); mem_filters(13)(149) <= to_signed(0,32); mem_filters(13)(150) <= to_signed(0,32);
  mem_filters(13)(151) <= to_signed(0,32); mem_filters(13)(152) <= to_signed(0,32); mem_filters(13)(153) <= to_signed(0,32);
  mem_filters(13)(154) <= to_signed(0,32); mem_filters(13)(155) <= to_signed(0,32); mem_filters(13)(156) <= to_signed(0,32);
  mem_filters(13)(157) <= to_signed(0,32); mem_filters(13)(158) <= to_signed(0,32); mem_filters(13)(159) <= to_signed(0,32);
  mem_filters(13)(160) <= to_signed(0,32); mem_filters(13)(161) <= to_signed(0,32); mem_filters(13)(162) <= to_signed(0,32);
  mem_filters(13)(163) <= to_signed(0,32); mem_filters(13)(164) <= to_signed(0,32); mem_filters(13)(165) <= to_signed(0,32);
  mem_filters(13)(166) <= to_signed(0,32); mem_filters(13)(167) <= to_signed(0,32); mem_filters(13)(168) <= to_signed(0,32);
  mem_filters(13)(169) <= to_signed(0,32); mem_filters(13)(170) <= to_signed(0,32); mem_filters(13)(171) <= to_signed(0,32);
  mem_filters(13)(172) <= to_signed(0,32); mem_filters(13)(173) <= to_signed(0,32); mem_filters(13)(174) <= to_signed(0,32);
  mem_filters(13)(175) <= to_signed(0,32); mem_filters(13)(176) <= to_signed(0,32); mem_filters(13)(177) <= to_signed(0,32);
  mem_filters(13)(178) <= to_signed(0,32); mem_filters(13)(179) <= to_signed(0,32); mem_filters(13)(180) <= to_signed(0,32);
  mem_filters(13)(181) <= to_signed(0,32); mem_filters(13)(182) <= to_signed(0,32); mem_filters(13)(183) <= to_signed(0,32);
  mem_filters(13)(184) <= to_signed(0,32); mem_filters(13)(185) <= to_signed(0,32); mem_filters(13)(186) <= to_signed(0,32);
  mem_filters(13)(187) <= to_signed(0,32); mem_filters(13)(188) <= to_signed(0,32); mem_filters(13)(189) <= to_signed(0,32);
  mem_filters(13)(190) <= to_signed(0,32); mem_filters(13)(191) <= to_signed(0,32); mem_filters(13)(192) <= to_signed(0,32);
  mem_filters(13)(193) <= to_signed(0,32); mem_filters(13)(194) <= to_signed(0,32); mem_filters(13)(195) <= to_signed(0,32);
  mem_filters(13)(196) <= to_signed(0,32); mem_filters(13)(197) <= to_signed(0,32); mem_filters(13)(198) <= to_signed(0,32);
  mem_filters(13)(199) <= to_signed(0,32); mem_filters(13)(200) <= to_signed(0,32); mem_filters(13)(201) <= to_signed(0,32);
  mem_filters(13)(202) <= to_signed(0,32); mem_filters(13)(203) <= to_signed(0,32); mem_filters(13)(204) <= to_signed(0,32);
  mem_filters(13)(205) <= to_signed(0,32); mem_filters(13)(206) <= to_signed(0,32); mem_filters(13)(207) <= to_signed(0,32);
  mem_filters(13)(208) <= to_signed(0,32); mem_filters(13)(209) <= to_signed(0,32); mem_filters(13)(210) <= to_signed(0,32);
  mem_filters(13)(211) <= to_signed(0,32); mem_filters(13)(212) <= to_signed(0,32); mem_filters(13)(213) <= to_signed(0,32);
  mem_filters(13)(214) <= to_signed(0,32); mem_filters(13)(215) <= to_signed(0,32); mem_filters(13)(216) <= to_signed(0,32);
  mem_filters(13)(217) <= to_signed(0,32); mem_filters(13)(218) <= to_signed(0,32); mem_filters(13)(219) <= to_signed(0,32);
  mem_filters(13)(220) <= to_signed(0,32); mem_filters(13)(221) <= to_signed(0,32); mem_filters(13)(222) <= to_signed(0,32);
  mem_filters(13)(223) <= to_signed(0,32); mem_filters(13)(224) <= to_signed(0,32); mem_filters(13)(225) <= to_signed(0,32);
  mem_filters(13)(226) <= to_signed(0,32); mem_filters(13)(227) <= to_signed(0,32); mem_filters(13)(228) <= to_signed(0,32);
  mem_filters(13)(229) <= to_signed(0,32); mem_filters(13)(230) <= to_signed(0,32); mem_filters(13)(231) <= to_signed(0,32);
  mem_filters(13)(232) <= to_signed(0,32); mem_filters(13)(233) <= to_signed(0,32); mem_filters(13)(234) <= to_signed(0,32);
  mem_filters(13)(235) <= to_signed(0,32); mem_filters(13)(236) <= to_signed(0,32); mem_filters(13)(237) <= to_signed(0,32);
  mem_filters(13)(238) <= to_signed(0,32); mem_filters(13)(239) <= to_signed(0,32); mem_filters(13)(240) <= to_signed(0,32);
  mem_filters(13)(241) <= to_signed(0,32); mem_filters(13)(242) <= to_signed(0,32); mem_filters(13)(243) <= to_signed(0,32);
  mem_filters(13)(244) <= to_signed(0,32); mem_filters(13)(245) <= to_signed(0,32); mem_filters(13)(246) <= to_signed(0,32);
  mem_filters(13)(247) <= to_signed(0,32); mem_filters(13)(248) <= to_signed(0,32); mem_filters(13)(249) <= to_signed(0,32);
  mem_filters(13)(250) <= to_signed(0,32); mem_filters(13)(251) <= to_signed(0,32); mem_filters(13)(252) <= to_signed(0,32);
  mem_filters(13)(253) <= to_signed(0,32); mem_filters(13)(254) <= to_signed(0,32); mem_filters(13)(255) <= to_signed(0,32);
  
  --Filter 14
  mem_filters(14)(0) <= to_signed(0,32); mem_filters(14)(1) <= to_signed(0,32); mem_filters(14)(2) <= to_signed(0,32);
  mem_filters(14)(3) <= to_signed(0,32); mem_filters(14)(4) <= to_signed(0,32); mem_filters(14)(5) <= to_signed(0,32);
  mem_filters(14)(6) <= to_signed(0,32); mem_filters(14)(7) <= to_signed(0,32); mem_filters(14)(8) <= to_signed(0,32);
  mem_filters(14)(9) <= to_signed(0,32); mem_filters(14)(10) <= to_signed(0,32); mem_filters(14)(11) <= to_signed(0,32);
  mem_filters(14)(12) <= to_signed(0,32); mem_filters(14)(13) <= to_signed(0,32); mem_filters(14)(14) <= to_signed(0,32);
  mem_filters(14)(15) <= to_signed(0,32); mem_filters(14)(16) <= to_signed(0,32); mem_filters(14)(17) <= to_signed(0,32);
  mem_filters(14)(18) <= to_signed(0,32); mem_filters(14)(19) <= to_signed(0,32); mem_filters(14)(20) <= to_signed(0,32);
  mem_filters(14)(21) <= to_signed(0,32); mem_filters(14)(22) <= to_signed(0,32); mem_filters(14)(23) <= to_signed(0,32);
  mem_filters(14)(24) <= to_signed(0,32); mem_filters(14)(25) <= to_signed(0,32); mem_filters(14)(26) <= to_signed(0,32);
  mem_filters(14)(27) <= to_signed(0,32); mem_filters(14)(28) <= to_signed(0,32); mem_filters(14)(29) <= to_signed(0,32);
  mem_filters(14)(30) <= to_signed(0,32); mem_filters(14)(31) <= to_signed(0,32); mem_filters(14)(32) <= to_signed(0,32);
  mem_filters(14)(33) <= to_signed(0,32); mem_filters(14)(34) <= to_signed(0,32); mem_filters(14)(35) <= to_signed(0,32);
  mem_filters(14)(36) <= to_signed(0,32); mem_filters(14)(37) <= to_signed(0,32); mem_filters(14)(38) <= to_signed(0,32);
  mem_filters(14)(39) <= to_signed(0,32); mem_filters(14)(40) <= to_signed(0,32); mem_filters(14)(41) <= to_signed(0,32);
  mem_filters(14)(42) <= to_signed(0,32); mem_filters(14)(43) <= to_signed(0,32); mem_filters(14)(44) <= to_signed(0,32);
  mem_filters(14)(45) <= to_signed(0,32);
  mem_filters(14)(46) <= to_signed(0,32); mem_filters(14)(47) <= to_signed(0,32); mem_filters(14)(48) <= to_signed(0,32);
  mem_filters(14)(49) <= to_signed(0,32); mem_filters(14)(50) <= to_signed(0,32); mem_filters(14)(51) <= to_signed(0,32);
  mem_filters(14)(52) <= to_signed(0,32); mem_filters(14)(53) <= to_signed(0,32); mem_filters(14)(54) <= to_signed(0,32);
  mem_filters(14)(55) <= to_signed(0,32); mem_filters(14)(56) <= to_signed(0,32); mem_filters(14)(57) <= to_signed(0,32);
  mem_filters(14)(58) <= to_signed(0,32); mem_filters(14)(59) <= to_signed(0,32); mem_filters(14)(60) <= to_signed(0,32);
  mem_filters(14)(61) <= to_signed(0,32); mem_filters(14)(62) <= to_signed(0,32); mem_filters(14)(63) <= to_signed(0,32);
  mem_filters(14)(64) <= to_signed(0,32); mem_filters(14)(65) <= to_signed(0,32); mem_filters(14)(66) <= to_signed(0,32);
  mem_filters(14)(67) <= to_signed(0,32); mem_filters(14)(68) <= to_signed(0,32); mem_filters(14)(69) <= to_signed(0,32);
  mem_filters(14)(70) <= to_signed(0,32); mem_filters(14)(71) <= to_signed(0,32); mem_filters(14)(72) <= to_signed(0,32);
  mem_filters(14)(73) <= to_signed(0,32); mem_filters(14)(74) <= to_signed(0,32); mem_filters(14)(75) <= to_signed(0,32);
  mem_filters(14)(76) <= to_signed(0,32); mem_filters(14)(77) <= to_signed(0,32); mem_filters(14)(78) <= to_signed(0,32);
  mem_filters(14)(79) <= to_signed(0,32); mem_filters(14)(80) <= to_signed(0,32); mem_filters(14)(81) <= to_signed(0,32);
  mem_filters(14)(82) <= to_signed(0,32); mem_filters(14)(83) <= to_signed(0,32); mem_filters(14)(84) <= to_signed(0,32);
  mem_filters(14)(85) <= to_signed(0,32); mem_filters(14)(86) <= to_signed(0,32); mem_filters(14)(87) <= to_signed(0,32);
  mem_filters(14)(88) <= to_signed(0,32); mem_filters(14)(89) <= to_signed(0,32); mem_filters(14)(90) <= to_signed(0,32);
  mem_filters(14)(91) <= to_signed(0,32); mem_filters(14)(92) <= to_signed(0,32); mem_filters(14)(93) <= to_signed(0,32);
  mem_filters(14)(94) <= to_signed(0,32); mem_filters(14)(95) <= to_signed(0,32); mem_filters(14)(96) <= to_signed(0,32);
  mem_filters(14)(97) <= to_signed(0,32); mem_filters(14)(98) <= to_signed(0,32); mem_filters(14)(99) <= to_signed(0,32);
  mem_filters(14)(100) <= to_signed(0,32); mem_filters(14)(101) <= to_signed(0,32); mem_filters(14)(102) <= to_signed(0,32);
  mem_filters(14)(103) <= to_signed(0,32); mem_filters(14)(104) <= to_signed(0,32); mem_filters(14)(105) <= to_signed(0,32);
  mem_filters(14)(106) <= to_signed(0,32); mem_filters(14)(107) <= to_signed(0,32); mem_filters(14)(108) <= to_signed(0,32);
  mem_filters(14)(109) <= to_signed(0,32); mem_filters(14)(110) <= to_signed(0,32); mem_filters(14)(111) <= to_signed(0,32);
  mem_filters(14)(112) <= to_signed(0,32); mem_filters(14)(113) <= to_signed(0,32); mem_filters(14)(114) <= to_signed(0,32);
  mem_filters(14)(115) <= to_signed(0,32); mem_filters(14)(116) <= to_signed(0,32); mem_filters(14)(117) <= to_signed(0,32);
  mem_filters(14)(118) <= to_signed(0,32); mem_filters(14)(119) <= to_signed(0,32); mem_filters(14)(120) <= to_signed(0,32);
  mem_filters(14)(121) <= to_signed(0,32); mem_filters(14)(122) <= to_signed(0,32); mem_filters(14)(123) <= to_signed(0,32);
  mem_filters(14)(124) <= to_signed(0,32); mem_filters(14)(125) <= to_signed(0,32); mem_filters(14)(126) <= to_signed(0,32);
  mem_filters(14)(127) <= to_signed(0,32); mem_filters(14)(128) <= to_signed(0,32); mem_filters(14)(129) <= to_signed(0,32);
  mem_filters(14)(130) <= to_signed(0,32); mem_filters(14)(131) <= to_signed(0,32); mem_filters(14)(132) <= to_signed(0,32);
  mem_filters(14)(133) <= to_signed(0,32); mem_filters(14)(134) <= to_signed(0,32); mem_filters(14)(135) <= to_signed(0,32);
  mem_filters(14)(136) <= to_signed(0,32); mem_filters(14)(137) <= to_signed(0,32); mem_filters(14)(138) <= to_signed(0,32);
  mem_filters(14)(139) <= to_signed(0,32); mem_filters(14)(140) <= to_signed(0,32); mem_filters(14)(141) <= to_signed(0,32);
  mem_filters(14)(142) <= to_signed(0,32); mem_filters(14)(143) <= to_signed(0,32); mem_filters(14)(144) <= to_signed(0,32);
  mem_filters(14)(145) <= to_signed(0,32); mem_filters(14)(146) <= to_signed(0,32); mem_filters(14)(147) <= to_signed(0,32);
  mem_filters(14)(148) <= to_signed(0,32); mem_filters(14)(149) <= to_signed(0,32); mem_filters(14)(150) <= to_signed(0,32);
  mem_filters(14)(151) <= to_signed(0,32); mem_filters(14)(152) <= to_signed(0,32); mem_filters(14)(153) <= to_signed(0,32);
  mem_filters(14)(154) <= to_signed(0,32); mem_filters(14)(155) <= to_signed(0,32); mem_filters(14)(156) <= to_signed(0,32);
  mem_filters(14)(157) <= to_signed(0,32); mem_filters(14)(158) <= to_signed(0,32); mem_filters(14)(159) <= to_signed(0,32);
  mem_filters(14)(160) <= to_signed(0,32); mem_filters(14)(161) <= to_signed(0,32); mem_filters(14)(162) <= to_signed(0,32);
  mem_filters(14)(163) <= to_signed(0,32); mem_filters(14)(164) <= to_signed(0,32); mem_filters(14)(165) <= to_signed(0,32);
  mem_filters(14)(166) <= to_signed(0,32); mem_filters(14)(167) <= to_signed(0,32); mem_filters(14)(168) <= to_signed(0,32);
  mem_filters(14)(169) <= to_signed(0,32); mem_filters(14)(170) <= to_signed(0,32); mem_filters(14)(171) <= to_signed(0,32);
  mem_filters(14)(172) <= to_signed(0,32); mem_filters(14)(173) <= to_signed(0,32); mem_filters(14)(174) <= to_signed(0,32);
  mem_filters(14)(175) <= to_signed(0,32); mem_filters(14)(176) <= to_signed(0,32); mem_filters(14)(177) <= to_signed(0,32);
  mem_filters(14)(178) <= to_signed(0,32); mem_filters(14)(179) <= to_signed(0,32); mem_filters(14)(180) <= to_signed(0,32);
  mem_filters(14)(181) <= to_signed(0,32); mem_filters(14)(182) <= to_signed(0,32); mem_filters(14)(183) <= to_signed(0,32);
  mem_filters(14)(184) <= to_signed(0,32); mem_filters(14)(185) <= to_signed(0,32); mem_filters(14)(186) <= to_signed(0,32);
  mem_filters(14)(187) <= to_signed(0,32); mem_filters(14)(188) <= to_signed(0,32); mem_filters(14)(189) <= to_signed(0,32);
  mem_filters(14)(190) <= to_signed(0,32); mem_filters(14)(191) <= to_signed(0,32); mem_filters(14)(192) <= to_signed(0,32);
  mem_filters(14)(193) <= to_signed(0,32); mem_filters(14)(194) <= to_signed(0,32); mem_filters(14)(195) <= to_signed(0,32);
  mem_filters(14)(196) <= to_signed(0,32); mem_filters(14)(197) <= to_signed(0,32); mem_filters(14)(198) <= to_signed(0,32);
  mem_filters(14)(199) <= to_signed(0,32); mem_filters(14)(200) <= to_signed(0,32); mem_filters(14)(201) <= to_signed(0,32);
  mem_filters(14)(202) <= to_signed(0,32); mem_filters(14)(203) <= to_signed(0,32); mem_filters(14)(204) <= to_signed(0,32);
  mem_filters(14)(205) <= to_signed(0,32); mem_filters(14)(206) <= to_signed(0,32); mem_filters(14)(207) <= to_signed(0,32);
  mem_filters(14)(208) <= to_signed(0,32); mem_filters(14)(209) <= to_signed(0,32); mem_filters(14)(210) <= to_signed(0,32);
  mem_filters(14)(211) <= to_signed(0,32); mem_filters(14)(212) <= to_signed(0,32); mem_filters(14)(213) <= to_signed(0,32);
  mem_filters(14)(214) <= to_signed(0,32); mem_filters(14)(215) <= to_signed(0,32); mem_filters(14)(216) <= to_signed(0,32);
  mem_filters(14)(217) <= to_signed(0,32); mem_filters(14)(218) <= to_signed(0,32); mem_filters(14)(219) <= to_signed(0,32);
  mem_filters(14)(220) <= to_signed(0,32); mem_filters(14)(221) <= to_signed(0,32); mem_filters(14)(222) <= to_signed(0,32);
  mem_filters(14)(223) <= to_signed(0,32); mem_filters(14)(224) <= to_signed(0,32); mem_filters(14)(225) <= to_signed(0,32);
  mem_filters(14)(226) <= to_signed(0,32); mem_filters(14)(227) <= to_signed(0,32); mem_filters(14)(228) <= to_signed(0,32);
  mem_filters(14)(229) <= to_signed(0,32); mem_filters(14)(230) <= to_signed(0,32); mem_filters(14)(231) <= to_signed(0,32);
  mem_filters(14)(232) <= to_signed(0,32); mem_filters(14)(233) <= to_signed(0,32); mem_filters(14)(234) <= to_signed(0,32);
  mem_filters(14)(235) <= to_signed(0,32); mem_filters(14)(236) <= to_signed(0,32); mem_filters(14)(237) <= to_signed(0,32);
  mem_filters(14)(238) <= to_signed(0,32); mem_filters(14)(239) <= to_signed(0,32); mem_filters(14)(240) <= to_signed(0,32);
  mem_filters(14)(241) <= to_signed(0,32); mem_filters(14)(242) <= to_signed(0,32); mem_filters(14)(243) <= to_signed(0,32);
  mem_filters(14)(244) <= to_signed(0,32); mem_filters(14)(245) <= to_signed(0,32); mem_filters(14)(246) <= to_signed(0,32);
  mem_filters(14)(247) <= to_signed(0,32); mem_filters(14)(248) <= to_signed(0,32); mem_filters(14)(249) <= to_signed(0,32);
  mem_filters(14)(250) <= to_signed(0,32); mem_filters(14)(251) <= to_signed(0,32); mem_filters(14)(252) <= to_signed(0,32);
  mem_filters(14)(253) <= to_signed(0,32); mem_filters(14)(254) <= to_signed(0,32); mem_filters(14)(255) <= to_signed(0,32);
  
  --Filter 15
  mem_filters(15)(0) <= to_signed(0,32); mem_filters(15)(1) <= to_signed(0,32); mem_filters(15)(2) <= to_signed(0,32);
  mem_filters(15)(3) <= to_signed(0,32); mem_filters(15)(4) <= to_signed(0,32); mem_filters(15)(5) <= to_signed(0,32);
  mem_filters(15)(6) <= to_signed(0,32); mem_filters(15)(7) <= to_signed(0,32); mem_filters(15)(8) <= to_signed(0,32);
  mem_filters(15)(9) <= to_signed(0,32); mem_filters(15)(10) <= to_signed(0,32); mem_filters(15)(11) <= to_signed(0,32);
  mem_filters(15)(12) <= to_signed(0,32); mem_filters(15)(13) <= to_signed(0,32); mem_filters(15)(14) <= to_signed(0,32);
  mem_filters(15)(15) <= to_signed(0,32); mem_filters(15)(16) <= to_signed(0,32); mem_filters(15)(17) <= to_signed(0,32);
  mem_filters(15)(18) <= to_signed(0,32); mem_filters(15)(19) <= to_signed(0,32); mem_filters(15)(20) <= to_signed(0,32);
  mem_filters(15)(21) <= to_signed(0,32); mem_filters(15)(22) <= to_signed(0,32); mem_filters(15)(23) <= to_signed(0,32);
  mem_filters(15)(24) <= to_signed(0,32); mem_filters(15)(25) <= to_signed(0,32); mem_filters(15)(26) <= to_signed(0,32);
  mem_filters(15)(27) <= to_signed(0,32); mem_filters(15)(28) <= to_signed(0,32); mem_filters(15)(29) <= to_signed(0,32);
  mem_filters(15)(30) <= to_signed(0,32); mem_filters(15)(31) <= to_signed(0,32); mem_filters(15)(32) <= to_signed(0,32);
  mem_filters(15)(33) <= to_signed(0,32); mem_filters(15)(34) <= to_signed(0,32); mem_filters(15)(35) <= to_signed(0,32);
  mem_filters(15)(36) <= to_signed(0,32); mem_filters(15)(37) <= to_signed(0,32); mem_filters(15)(38) <= to_signed(0,32);
  mem_filters(15)(39) <= to_signed(0,32); mem_filters(15)(40) <= to_signed(0,32); mem_filters(15)(41) <= to_signed(0,32);
  mem_filters(15)(42) <= to_signed(0,32); mem_filters(15)(43) <= to_signed(0,32); mem_filters(15)(44) <= to_signed(0,32);
  mem_filters(15)(45) <= to_signed(0,32);
  mem_filters(15)(46) <= to_signed(0,32); mem_filters(15)(47) <= to_signed(0,32); mem_filters(15)(48) <= to_signed(0,32);
  mem_filters(15)(49) <= to_signed(0,32); mem_filters(15)(50) <= to_signed(0,32); mem_filters(15)(51) <= to_signed(0,32);
  mem_filters(15)(52) <= to_signed(0,32); mem_filters(15)(53) <= to_signed(0,32); mem_filters(15)(54) <= to_signed(0,32);
  mem_filters(15)(55) <= to_signed(0,32); mem_filters(15)(56) <= to_signed(0,32); mem_filters(15)(57) <= to_signed(0,32);
  mem_filters(15)(58) <= to_signed(0,32); mem_filters(15)(59) <= to_signed(0,32); mem_filters(15)(60) <= to_signed(0,32);
  mem_filters(15)(61) <= to_signed(0,32); mem_filters(15)(62) <= to_signed(0,32); mem_filters(15)(63) <= to_signed(0,32);
  mem_filters(15)(64) <= to_signed(0,32); mem_filters(15)(65) <= to_signed(0,32); mem_filters(15)(66) <= to_signed(0,32);
  mem_filters(15)(67) <= to_signed(0,32); mem_filters(15)(68) <= to_signed(0,32); mem_filters(15)(69) <= to_signed(0,32);
  mem_filters(15)(70) <= to_signed(0,32); mem_filters(15)(71) <= to_signed(0,32); mem_filters(15)(72) <= to_signed(0,32);
  mem_filters(15)(73) <= to_signed(0,32); mem_filters(15)(74) <= to_signed(0,32); mem_filters(15)(75) <= to_signed(0,32);
  mem_filters(15)(76) <= to_signed(0,32); mem_filters(15)(77) <= to_signed(0,32); mem_filters(15)(78) <= to_signed(0,32);
  mem_filters(15)(79) <= to_signed(0,32); mem_filters(15)(80) <= to_signed(0,32); mem_filters(15)(81) <= to_signed(0,32);
  mem_filters(15)(82) <= to_signed(0,32); mem_filters(15)(83) <= to_signed(0,32); mem_filters(15)(84) <= to_signed(0,32);
  mem_filters(15)(85) <= to_signed(0,32); mem_filters(15)(86) <= to_signed(0,32); mem_filters(15)(87) <= to_signed(0,32);
  mem_filters(15)(88) <= to_signed(0,32); mem_filters(15)(89) <= to_signed(0,32); mem_filters(15)(90) <= to_signed(0,32);
  mem_filters(15)(91) <= to_signed(0,32); mem_filters(15)(92) <= to_signed(0,32); mem_filters(15)(93) <= to_signed(0,32);
  mem_filters(15)(94) <= to_signed(0,32); mem_filters(15)(95) <= to_signed(0,32); mem_filters(15)(96) <= to_signed(0,32);
  mem_filters(15)(97) <= to_signed(0,32); mem_filters(15)(98) <= to_signed(0,32); mem_filters(15)(99) <= to_signed(0,32);
  mem_filters(15)(100) <= to_signed(0,32); mem_filters(15)(101) <= to_signed(0,32); mem_filters(15)(102) <= to_signed(0,32);
  mem_filters(15)(103) <= to_signed(0,32); mem_filters(15)(104) <= to_signed(0,32); mem_filters(15)(105) <= to_signed(0,32);
  mem_filters(15)(106) <= to_signed(0,32); mem_filters(15)(107) <= to_signed(0,32); mem_filters(15)(108) <= to_signed(0,32);
  mem_filters(15)(109) <= to_signed(0,32); mem_filters(15)(110) <= to_signed(0,32); mem_filters(15)(111) <= to_signed(0,32);
  mem_filters(15)(112) <= to_signed(0,32); mem_filters(15)(113) <= to_signed(0,32); mem_filters(15)(114) <= to_signed(0,32);
  mem_filters(15)(115) <= to_signed(0,32); mem_filters(15)(116) <= to_signed(0,32); mem_filters(15)(117) <= to_signed(0,32);
  mem_filters(15)(118) <= to_signed(0,32); mem_filters(15)(119) <= to_signed(0,32); mem_filters(15)(120) <= to_signed(0,32);
  mem_filters(15)(121) <= to_signed(0,32); mem_filters(15)(122) <= to_signed(0,32); mem_filters(15)(123) <= to_signed(0,32);
  mem_filters(15)(124) <= to_signed(0,32); mem_filters(15)(125) <= to_signed(0,32); mem_filters(15)(126) <= to_signed(0,32);
  mem_filters(15)(127) <= to_signed(0,32); mem_filters(15)(128) <= to_signed(0,32); mem_filters(15)(129) <= to_signed(0,32);
  mem_filters(15)(130) <= to_signed(0,32); mem_filters(15)(131) <= to_signed(0,32); mem_filters(15)(132) <= to_signed(0,32);
  mem_filters(15)(133) <= to_signed(0,32); mem_filters(15)(134) <= to_signed(0,32); mem_filters(15)(135) <= to_signed(0,32);
  mem_filters(15)(136) <= to_signed(0,32); mem_filters(15)(137) <= to_signed(0,32); mem_filters(15)(138) <= to_signed(0,32);
  mem_filters(15)(139) <= to_signed(0,32); mem_filters(15)(140) <= to_signed(0,32); mem_filters(15)(141) <= to_signed(0,32);
  mem_filters(15)(142) <= to_signed(0,32); mem_filters(15)(143) <= to_signed(0,32); mem_filters(15)(144) <= to_signed(0,32);
  mem_filters(15)(145) <= to_signed(0,32); mem_filters(15)(146) <= to_signed(0,32); mem_filters(15)(147) <= to_signed(0,32);
  mem_filters(15)(148) <= to_signed(0,32); mem_filters(15)(149) <= to_signed(0,32); mem_filters(15)(150) <= to_signed(0,32);
  mem_filters(15)(151) <= to_signed(0,32); mem_filters(15)(152) <= to_signed(0,32); mem_filters(15)(153) <= to_signed(0,32);
  mem_filters(15)(154) <= to_signed(0,32); mem_filters(15)(155) <= to_signed(0,32); mem_filters(15)(156) <= to_signed(0,32);
  mem_filters(15)(157) <= to_signed(0,32); mem_filters(15)(158) <= to_signed(0,32); mem_filters(15)(159) <= to_signed(0,32);
  mem_filters(15)(160) <= to_signed(0,32); mem_filters(15)(161) <= to_signed(0,32); mem_filters(15)(162) <= to_signed(0,32);
  mem_filters(15)(163) <= to_signed(0,32); mem_filters(15)(164) <= to_signed(0,32); mem_filters(15)(165) <= to_signed(0,32);
  mem_filters(15)(166) <= to_signed(0,32); mem_filters(15)(167) <= to_signed(0,32); mem_filters(15)(168) <= to_signed(0,32);
  mem_filters(15)(169) <= to_signed(0,32); mem_filters(15)(170) <= to_signed(0,32); mem_filters(15)(171) <= to_signed(0,32);
  mem_filters(15)(172) <= to_signed(0,32); mem_filters(15)(173) <= to_signed(0,32); mem_filters(15)(174) <= to_signed(0,32);
  mem_filters(15)(175) <= to_signed(0,32); mem_filters(15)(176) <= to_signed(0,32); mem_filters(15)(177) <= to_signed(0,32);
  mem_filters(15)(178) <= to_signed(0,32); mem_filters(15)(179) <= to_signed(0,32); mem_filters(15)(180) <= to_signed(0,32);
  mem_filters(15)(181) <= to_signed(0,32); mem_filters(15)(182) <= to_signed(0,32); mem_filters(15)(183) <= to_signed(0,32);
  mem_filters(15)(184) <= to_signed(0,32); mem_filters(15)(185) <= to_signed(0,32); mem_filters(15)(186) <= to_signed(0,32);
  mem_filters(15)(187) <= to_signed(0,32); mem_filters(15)(188) <= to_signed(0,32); mem_filters(15)(189) <= to_signed(0,32);
  mem_filters(15)(190) <= to_signed(0,32); mem_filters(15)(191) <= to_signed(0,32); mem_filters(15)(192) <= to_signed(0,32);
  mem_filters(15)(193) <= to_signed(0,32); mem_filters(15)(194) <= to_signed(0,32); mem_filters(15)(195) <= to_signed(0,32);
  mem_filters(15)(196) <= to_signed(0,32); mem_filters(15)(197) <= to_signed(0,32); mem_filters(15)(198) <= to_signed(0,32);
  mem_filters(15)(199) <= to_signed(0,32); mem_filters(15)(200) <= to_signed(0,32); mem_filters(15)(201) <= to_signed(0,32);
  mem_filters(15)(202) <= to_signed(0,32); mem_filters(15)(203) <= to_signed(0,32); mem_filters(15)(204) <= to_signed(0,32);
  mem_filters(15)(205) <= to_signed(0,32); mem_filters(15)(206) <= to_signed(0,32); mem_filters(15)(207) <= to_signed(0,32);
  mem_filters(15)(208) <= to_signed(0,32); mem_filters(15)(209) <= to_signed(0,32); mem_filters(15)(210) <= to_signed(0,32);
  mem_filters(15)(211) <= to_signed(0,32); mem_filters(15)(212) <= to_signed(0,32); mem_filters(15)(213) <= to_signed(0,32);
  mem_filters(15)(214) <= to_signed(0,32); mem_filters(15)(215) <= to_signed(0,32); mem_filters(15)(216) <= to_signed(0,32);
  mem_filters(15)(217) <= to_signed(0,32); mem_filters(15)(218) <= to_signed(0,32); mem_filters(15)(219) <= to_signed(0,32);
  mem_filters(15)(220) <= to_signed(0,32); mem_filters(15)(221) <= to_signed(0,32); mem_filters(15)(222) <= to_signed(0,32);
  mem_filters(15)(223) <= to_signed(0,32); mem_filters(15)(224) <= to_signed(0,32); mem_filters(15)(225) <= to_signed(0,32);
  mem_filters(15)(226) <= to_signed(0,32); mem_filters(15)(227) <= to_signed(0,32); mem_filters(15)(228) <= to_signed(0,32);
  mem_filters(15)(229) <= to_signed(0,32); mem_filters(15)(230) <= to_signed(0,32); mem_filters(15)(231) <= to_signed(0,32);
  mem_filters(15)(232) <= to_signed(0,32); mem_filters(15)(233) <= to_signed(0,32); mem_filters(15)(234) <= to_signed(0,32);
  mem_filters(15)(235) <= to_signed(0,32); mem_filters(15)(236) <= to_signed(0,32); mem_filters(15)(237) <= to_signed(0,32);
  mem_filters(15)(238) <= to_signed(0,32); mem_filters(15)(239) <= to_signed(0,32); mem_filters(15)(240) <= to_signed(0,32);
  mem_filters(15)(241) <= to_signed(0,32); mem_filters(15)(242) <= to_signed(0,32); mem_filters(15)(243) <= to_signed(0,32);
  mem_filters(15)(244) <= to_signed(0,32); mem_filters(15)(245) <= to_signed(0,32); mem_filters(15)(246) <= to_signed(0,32);
  mem_filters(15)(247) <= to_signed(0,32); mem_filters(15)(248) <= to_signed(0,32); mem_filters(15)(249) <= to_signed(0,32);
  mem_filters(15)(250) <= to_signed(0,32); mem_filters(15)(251) <= to_signed(0,32); mem_filters(15)(252) <= to_signed(0,32);
  mem_filters(15)(253) <= to_signed(0,32); mem_filters(15)(254) <= to_signed(0,32); mem_filters(15)(255) <= to_signed(0,32);
  
  --Filter 16
  mem_filters(16)(0) <= to_signed(0,32); mem_filters(16)(1) <= to_signed(0,32); mem_filters(16)(2) <= to_signed(0,32);
  mem_filters(16)(3) <= to_signed(0,32); mem_filters(16)(4) <= to_signed(0,32); mem_filters(16)(5) <= to_signed(0,32);
  mem_filters(16)(6) <= to_signed(0,32); mem_filters(16)(7) <= to_signed(0,32); mem_filters(16)(8) <= to_signed(0,32);
  mem_filters(16)(9) <= to_signed(0,32); mem_filters(16)(10) <= to_signed(0,32); mem_filters(16)(11) <= to_signed(0,32);
  mem_filters(16)(12) <= to_signed(0,32); mem_filters(16)(13) <= to_signed(0,32); mem_filters(16)(14) <= to_signed(0,32);
  mem_filters(16)(15) <= to_signed(0,32); mem_filters(16)(16) <= to_signed(0,32); mem_filters(16)(17) <= to_signed(0,32);
  mem_filters(16)(18) <= to_signed(0,32); mem_filters(16)(19) <= to_signed(0,32); mem_filters(16)(20) <= to_signed(0,32);
  mem_filters(16)(21) <= to_signed(0,32); mem_filters(16)(22) <= to_signed(0,32); mem_filters(16)(23) <= to_signed(0,32);
  mem_filters(16)(24) <= to_signed(0,32); mem_filters(16)(25) <= to_signed(0,32); mem_filters(16)(26) <= to_signed(0,32);
  mem_filters(16)(27) <= to_signed(0,32); mem_filters(16)(28) <= to_signed(0,32); mem_filters(16)(29) <= to_signed(0,32);
  mem_filters(16)(30) <= to_signed(0,32); mem_filters(16)(31) <= to_signed(0,32); mem_filters(16)(32) <= to_signed(0,32);
  mem_filters(16)(33) <= to_signed(0,32); mem_filters(16)(34) <= to_signed(0,32); mem_filters(16)(35) <= to_signed(0,32);
  mem_filters(16)(36) <= to_signed(0,32); mem_filters(16)(37) <= to_signed(0,32); mem_filters(16)(38) <= to_signed(0,32);
  mem_filters(16)(39) <= to_signed(0,32); mem_filters(16)(40) <= to_signed(0,32); mem_filters(16)(41) <= to_signed(0,32);
  mem_filters(16)(42) <= to_signed(0,32); mem_filters(16)(43) <= to_signed(0,32); mem_filters(16)(44) <= to_signed(0,32);
  mem_filters(16)(45) <= to_signed(0,32);
  mem_filters(16)(46) <= to_signed(0,32); mem_filters(16)(47) <= to_signed(0,32); mem_filters(16)(48) <= to_signed(0,32);
  mem_filters(16)(49) <= to_signed(0,32); mem_filters(16)(50) <= to_signed(0,32); mem_filters(16)(51) <= to_signed(0,32);
  mem_filters(16)(52) <= to_signed(0,32); mem_filters(16)(53) <= to_signed(0,32); mem_filters(16)(54) <= to_signed(0,32);
  mem_filters(16)(55) <= to_signed(0,32); mem_filters(16)(56) <= to_signed(0,32); mem_filters(16)(57) <= to_signed(0,32);
  mem_filters(16)(58) <= to_signed(0,32); mem_filters(16)(59) <= to_signed(0,32); mem_filters(16)(60) <= to_signed(0,32);
  mem_filters(16)(61) <= to_signed(0,32); mem_filters(16)(62) <= to_signed(0,32); mem_filters(16)(63) <= to_signed(0,32);
  mem_filters(16)(64) <= to_signed(0,32); mem_filters(16)(65) <= to_signed(0,32); mem_filters(16)(66) <= to_signed(0,32);
  mem_filters(16)(67) <= to_signed(0,32); mem_filters(16)(68) <= to_signed(0,32); mem_filters(16)(69) <= to_signed(0,32);
  mem_filters(16)(70) <= to_signed(0,32); mem_filters(16)(71) <= to_signed(0,32); mem_filters(16)(72) <= to_signed(0,32);
  mem_filters(16)(73) <= to_signed(0,32); mem_filters(16)(74) <= to_signed(0,32); mem_filters(16)(75) <= to_signed(0,32);
  mem_filters(16)(76) <= to_signed(0,32); mem_filters(16)(77) <= to_signed(0,32); mem_filters(16)(78) <= to_signed(0,32);
  mem_filters(16)(79) <= to_signed(0,32); mem_filters(16)(80) <= to_signed(0,32); mem_filters(16)(81) <= to_signed(0,32);
  mem_filters(16)(82) <= to_signed(0,32); mem_filters(16)(83) <= to_signed(0,32); mem_filters(16)(84) <= to_signed(0,32);
  mem_filters(16)(85) <= to_signed(0,32); mem_filters(16)(86) <= to_signed(0,32); mem_filters(16)(87) <= to_signed(0,32);
  mem_filters(16)(88) <= to_signed(0,32); mem_filters(16)(89) <= to_signed(0,32); mem_filters(16)(90) <= to_signed(0,32);
  mem_filters(16)(91) <= to_signed(0,32); mem_filters(16)(92) <= to_signed(0,32); mem_filters(16)(93) <= to_signed(0,32);
  mem_filters(16)(94) <= to_signed(0,32); mem_filters(16)(95) <= to_signed(0,32); mem_filters(16)(96) <= to_signed(0,32);
  mem_filters(16)(97) <= to_signed(0,32); mem_filters(16)(98) <= to_signed(0,32); mem_filters(16)(99) <= to_signed(0,32);
  mem_filters(16)(100) <= to_signed(0,32); mem_filters(16)(101) <= to_signed(0,32); mem_filters(16)(102) <= to_signed(0,32);
  mem_filters(16)(103) <= to_signed(0,32); mem_filters(16)(104) <= to_signed(0,32); mem_filters(16)(105) <= to_signed(0,32);
  mem_filters(16)(106) <= to_signed(0,32); mem_filters(16)(107) <= to_signed(0,32); mem_filters(16)(108) <= to_signed(0,32);
  mem_filters(16)(109) <= to_signed(0,32); mem_filters(16)(110) <= to_signed(0,32); mem_filters(16)(111) <= to_signed(0,32);
  mem_filters(16)(112) <= to_signed(0,32); mem_filters(16)(113) <= to_signed(0,32); mem_filters(16)(114) <= to_signed(0,32);
  mem_filters(16)(115) <= to_signed(0,32); mem_filters(16)(116) <= to_signed(0,32); mem_filters(16)(117) <= to_signed(0,32);
  mem_filters(16)(118) <= to_signed(0,32); mem_filters(16)(119) <= to_signed(0,32); mem_filters(16)(120) <= to_signed(0,32);
  mem_filters(16)(121) <= to_signed(0,32); mem_filters(16)(122) <= to_signed(0,32); mem_filters(16)(123) <= to_signed(0,32);
  mem_filters(16)(124) <= to_signed(0,32); mem_filters(16)(125) <= to_signed(0,32); mem_filters(16)(126) <= to_signed(0,32);
  mem_filters(16)(127) <= to_signed(0,32); mem_filters(16)(128) <= to_signed(0,32); mem_filters(16)(129) <= to_signed(0,32);
  mem_filters(16)(130) <= to_signed(0,32); mem_filters(16)(131) <= to_signed(0,32); mem_filters(16)(132) <= to_signed(0,32);
  mem_filters(16)(133) <= to_signed(0,32); mem_filters(16)(134) <= to_signed(0,32); mem_filters(16)(135) <= to_signed(0,32);
  mem_filters(16)(136) <= to_signed(0,32); mem_filters(16)(137) <= to_signed(0,32); mem_filters(16)(138) <= to_signed(0,32);
  mem_filters(16)(139) <= to_signed(0,32); mem_filters(16)(140) <= to_signed(0,32); mem_filters(16)(141) <= to_signed(0,32);
  mem_filters(16)(142) <= to_signed(0,32); mem_filters(16)(143) <= to_signed(0,32); mem_filters(16)(144) <= to_signed(0,32);
  mem_filters(16)(145) <= to_signed(0,32); mem_filters(16)(146) <= to_signed(0,32); mem_filters(16)(147) <= to_signed(0,32);
  mem_filters(16)(148) <= to_signed(0,32); mem_filters(16)(149) <= to_signed(0,32); mem_filters(16)(150) <= to_signed(0,32);
  mem_filters(16)(151) <= to_signed(0,32); mem_filters(16)(152) <= to_signed(0,32); mem_filters(16)(153) <= to_signed(0,32);
  mem_filters(16)(154) <= to_signed(0,32); mem_filters(16)(155) <= to_signed(0,32); mem_filters(16)(156) <= to_signed(0,32);
  mem_filters(16)(157) <= to_signed(0,32); mem_filters(16)(158) <= to_signed(0,32); mem_filters(16)(159) <= to_signed(0,32);
  mem_filters(16)(160) <= to_signed(0,32); mem_filters(16)(161) <= to_signed(0,32); mem_filters(16)(162) <= to_signed(0,32);
  mem_filters(16)(163) <= to_signed(0,32); mem_filters(16)(164) <= to_signed(0,32); mem_filters(16)(165) <= to_signed(0,32);
  mem_filters(16)(166) <= to_signed(0,32); mem_filters(16)(167) <= to_signed(0,32); mem_filters(16)(168) <= to_signed(0,32);
  mem_filters(16)(169) <= to_signed(0,32); mem_filters(16)(170) <= to_signed(0,32); mem_filters(16)(171) <= to_signed(0,32);
  mem_filters(16)(172) <= to_signed(0,32); mem_filters(16)(173) <= to_signed(0,32); mem_filters(16)(174) <= to_signed(0,32);
  mem_filters(16)(175) <= to_signed(0,32); mem_filters(16)(176) <= to_signed(0,32); mem_filters(16)(177) <= to_signed(0,32);
  mem_filters(16)(178) <= to_signed(0,32); mem_filters(16)(179) <= to_signed(0,32); mem_filters(16)(180) <= to_signed(0,32);
  mem_filters(16)(181) <= to_signed(0,32); mem_filters(16)(182) <= to_signed(0,32); mem_filters(16)(183) <= to_signed(0,32);
  mem_filters(16)(184) <= to_signed(0,32); mem_filters(16)(185) <= to_signed(0,32); mem_filters(16)(186) <= to_signed(0,32);
  mem_filters(16)(187) <= to_signed(0,32); mem_filters(16)(188) <= to_signed(0,32); mem_filters(16)(189) <= to_signed(0,32);
  mem_filters(16)(190) <= to_signed(0,32); mem_filters(16)(191) <= to_signed(0,32); mem_filters(16)(192) <= to_signed(0,32);
  mem_filters(16)(193) <= to_signed(0,32); mem_filters(16)(194) <= to_signed(0,32); mem_filters(16)(195) <= to_signed(0,32);
  mem_filters(16)(196) <= to_signed(0,32); mem_filters(16)(197) <= to_signed(0,32); mem_filters(16)(198) <= to_signed(0,32);
  mem_filters(16)(199) <= to_signed(0,32); mem_filters(16)(200) <= to_signed(0,32); mem_filters(16)(201) <= to_signed(0,32);
  mem_filters(16)(202) <= to_signed(0,32); mem_filters(16)(203) <= to_signed(0,32); mem_filters(16)(204) <= to_signed(0,32);
  mem_filters(16)(205) <= to_signed(0,32); mem_filters(16)(206) <= to_signed(0,32); mem_filters(16)(207) <= to_signed(0,32);
  mem_filters(16)(208) <= to_signed(0,32); mem_filters(16)(209) <= to_signed(0,32); mem_filters(16)(210) <= to_signed(0,32);
  mem_filters(16)(211) <= to_signed(0,32); mem_filters(16)(212) <= to_signed(0,32); mem_filters(16)(213) <= to_signed(0,32);
  mem_filters(16)(214) <= to_signed(0,32); mem_filters(16)(215) <= to_signed(0,32); mem_filters(16)(216) <= to_signed(0,32);
  mem_filters(16)(217) <= to_signed(0,32); mem_filters(16)(218) <= to_signed(0,32); mem_filters(16)(219) <= to_signed(0,32);
  mem_filters(16)(220) <= to_signed(0,32); mem_filters(16)(221) <= to_signed(0,32); mem_filters(16)(222) <= to_signed(0,32);
  mem_filters(16)(223) <= to_signed(0,32); mem_filters(16)(224) <= to_signed(0,32); mem_filters(16)(225) <= to_signed(0,32);
  mem_filters(16)(226) <= to_signed(0,32); mem_filters(16)(227) <= to_signed(0,32); mem_filters(16)(228) <= to_signed(0,32);
  mem_filters(16)(229) <= to_signed(0,32); mem_filters(16)(230) <= to_signed(0,32); mem_filters(16)(231) <= to_signed(0,32);
  mem_filters(16)(232) <= to_signed(0,32); mem_filters(16)(233) <= to_signed(0,32); mem_filters(16)(234) <= to_signed(0,32);
  mem_filters(16)(235) <= to_signed(0,32); mem_filters(16)(236) <= to_signed(0,32); mem_filters(16)(237) <= to_signed(0,32);
  mem_filters(16)(238) <= to_signed(0,32); mem_filters(16)(239) <= to_signed(0,32); mem_filters(16)(240) <= to_signed(0,32);
  mem_filters(16)(241) <= to_signed(0,32); mem_filters(16)(242) <= to_signed(0,32); mem_filters(16)(243) <= to_signed(0,32);
  mem_filters(16)(244) <= to_signed(0,32); mem_filters(16)(245) <= to_signed(0,32); mem_filters(16)(246) <= to_signed(0,32);
  mem_filters(16)(247) <= to_signed(0,32); mem_filters(16)(248) <= to_signed(0,32); mem_filters(16)(249) <= to_signed(0,32);
  mem_filters(16)(250) <= to_signed(0,32); mem_filters(16)(251) <= to_signed(0,32); mem_filters(16)(252) <= to_signed(0,32);
  mem_filters(16)(253) <= to_signed(0,32); mem_filters(16)(254) <= to_signed(0,32); mem_filters(16)(255) <= to_signed(0,32);
  
  --Filter 17
  mem_filters(17)(0) <= to_signed(0,32); mem_filters(17)(1) <= to_signed(0,32); mem_filters(17)(2) <= to_signed(0,32);
  mem_filters(17)(3) <= to_signed(0,32); mem_filters(17)(4) <= to_signed(0,32); mem_filters(17)(5) <= to_signed(0,32);
  mem_filters(17)(6) <= to_signed(0,32); mem_filters(17)(7) <= to_signed(0,32); mem_filters(17)(8) <= to_signed(0,32);
  mem_filters(17)(9) <= to_signed(0,32); mem_filters(17)(10) <= to_signed(0,32); mem_filters(17)(11) <= to_signed(0,32);
  mem_filters(17)(12) <= to_signed(0,32); mem_filters(17)(13) <= to_signed(0,32); mem_filters(17)(14) <= to_signed(0,32);
  mem_filters(17)(15) <= to_signed(0,32); mem_filters(17)(16) <= to_signed(0,32); mem_filters(17)(17) <= to_signed(0,32);
  mem_filters(17)(18) <= to_signed(0,32); mem_filters(17)(19) <= to_signed(0,32); mem_filters(17)(20) <= to_signed(0,32);
  mem_filters(17)(21) <= to_signed(0,32); mem_filters(17)(22) <= to_signed(0,32); mem_filters(17)(23) <= to_signed(0,32);
  mem_filters(17)(24) <= to_signed(0,32); mem_filters(17)(25) <= to_signed(0,32); mem_filters(17)(26) <= to_signed(0,32);
  mem_filters(17)(27) <= to_signed(0,32); mem_filters(17)(28) <= to_signed(0,32); mem_filters(17)(29) <= to_signed(0,32);
  mem_filters(17)(30) <= to_signed(0,32); mem_filters(17)(31) <= to_signed(0,32); mem_filters(17)(32) <= to_signed(0,32);
  mem_filters(17)(33) <= to_signed(0,32); mem_filters(17)(34) <= to_signed(0,32); mem_filters(17)(35) <= to_signed(0,32);
  mem_filters(17)(36) <= to_signed(0,32); mem_filters(17)(37) <= to_signed(0,32); mem_filters(17)(38) <= to_signed(0,32);
  mem_filters(17)(39) <= to_signed(0,32); mem_filters(17)(40) <= to_signed(0,32); mem_filters(17)(41) <= to_signed(0,32);
  mem_filters(17)(42) <= to_signed(0,32); mem_filters(17)(43) <= to_signed(0,32); mem_filters(17)(44) <= to_signed(0,32);
  mem_filters(17)(45) <= to_signed(0,32);
  mem_filters(17)(46) <= to_signed(0,32); mem_filters(17)(47) <= to_signed(0,32); mem_filters(17)(48) <= to_signed(0,32);
  mem_filters(17)(49) <= to_signed(0,32); mem_filters(17)(50) <= to_signed(0,32); mem_filters(17)(51) <= to_signed(0,32);
  mem_filters(17)(52) <= to_signed(0,32); mem_filters(17)(53) <= to_signed(0,32); mem_filters(17)(54) <= to_signed(0,32);
  mem_filters(17)(55) <= to_signed(0,32); mem_filters(17)(56) <= to_signed(0,32); mem_filters(17)(57) <= to_signed(0,32);
  mem_filters(17)(58) <= to_signed(0,32); mem_filters(17)(59) <= to_signed(0,32); mem_filters(17)(60) <= to_signed(0,32);
  mem_filters(17)(61) <= to_signed(0,32); mem_filters(17)(62) <= to_signed(0,32); mem_filters(17)(63) <= to_signed(0,32);
  mem_filters(17)(64) <= to_signed(0,32); mem_filters(17)(65) <= to_signed(0,32); mem_filters(17)(66) <= to_signed(0,32);
  mem_filters(17)(67) <= to_signed(0,32); mem_filters(17)(68) <= to_signed(0,32); mem_filters(17)(69) <= to_signed(0,32);
  mem_filters(17)(70) <= to_signed(0,32); mem_filters(17)(71) <= to_signed(0,32); mem_filters(17)(72) <= to_signed(0,32);
  mem_filters(17)(73) <= to_signed(0,32); mem_filters(17)(74) <= to_signed(0,32); mem_filters(17)(75) <= to_signed(0,32);
  mem_filters(17)(76) <= to_signed(0,32); mem_filters(17)(77) <= to_signed(0,32); mem_filters(17)(78) <= to_signed(0,32);
  mem_filters(17)(79) <= to_signed(0,32); mem_filters(17)(80) <= to_signed(0,32); mem_filters(17)(81) <= to_signed(0,32);
  mem_filters(17)(82) <= to_signed(0,32); mem_filters(17)(83) <= to_signed(0,32); mem_filters(17)(84) <= to_signed(0,32);
  mem_filters(17)(85) <= to_signed(0,32); mem_filters(17)(86) <= to_signed(0,32); mem_filters(17)(87) <= to_signed(0,32);
  mem_filters(17)(88) <= to_signed(0,32); mem_filters(17)(89) <= to_signed(0,32); mem_filters(17)(90) <= to_signed(0,32);
  mem_filters(17)(91) <= to_signed(0,32); mem_filters(17)(92) <= to_signed(0,32); mem_filters(17)(93) <= to_signed(0,32);
  mem_filters(17)(94) <= to_signed(0,32); mem_filters(17)(95) <= to_signed(0,32); mem_filters(17)(96) <= to_signed(0,32);
  mem_filters(17)(97) <= to_signed(0,32); mem_filters(17)(98) <= to_signed(0,32); mem_filters(17)(99) <= to_signed(0,32);
  mem_filters(17)(100) <= to_signed(0,32); mem_filters(17)(101) <= to_signed(0,32); mem_filters(17)(102) <= to_signed(0,32);
  mem_filters(17)(103) <= to_signed(0,32); mem_filters(17)(104) <= to_signed(0,32); mem_filters(17)(105) <= to_signed(0,32);
  mem_filters(17)(106) <= to_signed(0,32); mem_filters(17)(107) <= to_signed(0,32); mem_filters(17)(108) <= to_signed(0,32);
  mem_filters(17)(109) <= to_signed(0,32); mem_filters(17)(110) <= to_signed(0,32); mem_filters(17)(111) <= to_signed(0,32);
  mem_filters(17)(112) <= to_signed(0,32); mem_filters(17)(113) <= to_signed(0,32); mem_filters(17)(114) <= to_signed(0,32);
  mem_filters(17)(115) <= to_signed(0,32); mem_filters(17)(116) <= to_signed(0,32); mem_filters(17)(117) <= to_signed(0,32);
  mem_filters(17)(118) <= to_signed(0,32); mem_filters(17)(119) <= to_signed(0,32); mem_filters(17)(120) <= to_signed(0,32);
  mem_filters(17)(121) <= to_signed(0,32); mem_filters(17)(122) <= to_signed(0,32); mem_filters(17)(123) <= to_signed(0,32);
  mem_filters(17)(124) <= to_signed(0,32); mem_filters(17)(125) <= to_signed(0,32); mem_filters(17)(126) <= to_signed(0,32);
  mem_filters(17)(127) <= to_signed(0,32); mem_filters(17)(128) <= to_signed(0,32); mem_filters(17)(129) <= to_signed(0,32);
  mem_filters(17)(130) <= to_signed(0,32); mem_filters(17)(131) <= to_signed(0,32); mem_filters(17)(132) <= to_signed(0,32);
  mem_filters(17)(133) <= to_signed(0,32); mem_filters(17)(134) <= to_signed(0,32); mem_filters(17)(135) <= to_signed(0,32);
  mem_filters(17)(136) <= to_signed(0,32); mem_filters(17)(137) <= to_signed(0,32); mem_filters(17)(138) <= to_signed(0,32);
  mem_filters(17)(139) <= to_signed(0,32); mem_filters(17)(140) <= to_signed(0,32); mem_filters(17)(141) <= to_signed(0,32);
  mem_filters(17)(142) <= to_signed(0,32); mem_filters(17)(143) <= to_signed(0,32); mem_filters(17)(144) <= to_signed(0,32);
  mem_filters(17)(145) <= to_signed(0,32); mem_filters(17)(146) <= to_signed(0,32); mem_filters(17)(147) <= to_signed(0,32);
  mem_filters(17)(148) <= to_signed(0,32); mem_filters(17)(149) <= to_signed(0,32); mem_filters(17)(150) <= to_signed(0,32);
  mem_filters(17)(151) <= to_signed(0,32); mem_filters(17)(152) <= to_signed(0,32); mem_filters(17)(153) <= to_signed(0,32);
  mem_filters(17)(154) <= to_signed(0,32); mem_filters(17)(155) <= to_signed(0,32); mem_filters(17)(156) <= to_signed(0,32);
  mem_filters(17)(157) <= to_signed(0,32); mem_filters(17)(158) <= to_signed(0,32); mem_filters(17)(159) <= to_signed(0,32);
  mem_filters(17)(160) <= to_signed(0,32); mem_filters(17)(161) <= to_signed(0,32); mem_filters(17)(162) <= to_signed(0,32);
  mem_filters(17)(163) <= to_signed(0,32); mem_filters(17)(164) <= to_signed(0,32); mem_filters(17)(165) <= to_signed(0,32);
  mem_filters(17)(166) <= to_signed(0,32); mem_filters(17)(167) <= to_signed(0,32); mem_filters(17)(168) <= to_signed(0,32);
  mem_filters(17)(169) <= to_signed(0,32); mem_filters(17)(170) <= to_signed(0,32); mem_filters(17)(171) <= to_signed(0,32);
  mem_filters(17)(172) <= to_signed(0,32); mem_filters(17)(173) <= to_signed(0,32); mem_filters(17)(174) <= to_signed(0,32);
  mem_filters(17)(175) <= to_signed(0,32); mem_filters(17)(176) <= to_signed(0,32); mem_filters(17)(177) <= to_signed(0,32);
  mem_filters(17)(178) <= to_signed(0,32); mem_filters(17)(179) <= to_signed(0,32); mem_filters(17)(180) <= to_signed(0,32);
  mem_filters(17)(181) <= to_signed(0,32); mem_filters(17)(182) <= to_signed(0,32); mem_filters(17)(183) <= to_signed(0,32);
  mem_filters(17)(184) <= to_signed(0,32); mem_filters(17)(185) <= to_signed(0,32); mem_filters(17)(186) <= to_signed(0,32);
  mem_filters(17)(187) <= to_signed(0,32); mem_filters(17)(188) <= to_signed(0,32); mem_filters(17)(189) <= to_signed(0,32);
  mem_filters(17)(190) <= to_signed(0,32); mem_filters(17)(191) <= to_signed(0,32); mem_filters(17)(192) <= to_signed(0,32);
  mem_filters(17)(193) <= to_signed(0,32); mem_filters(17)(194) <= to_signed(0,32); mem_filters(17)(195) <= to_signed(0,32);
  mem_filters(17)(196) <= to_signed(0,32); mem_filters(17)(197) <= to_signed(0,32); mem_filters(17)(198) <= to_signed(0,32);
  mem_filters(17)(199) <= to_signed(0,32); mem_filters(17)(200) <= to_signed(0,32); mem_filters(17)(201) <= to_signed(0,32);
  mem_filters(17)(202) <= to_signed(0,32); mem_filters(17)(203) <= to_signed(0,32); mem_filters(17)(204) <= to_signed(0,32);
  mem_filters(17)(205) <= to_signed(0,32); mem_filters(17)(206) <= to_signed(0,32); mem_filters(17)(207) <= to_signed(0,32);
  mem_filters(17)(208) <= to_signed(0,32); mem_filters(17)(209) <= to_signed(0,32); mem_filters(17)(210) <= to_signed(0,32);
  mem_filters(17)(211) <= to_signed(0,32); mem_filters(17)(212) <= to_signed(0,32); mem_filters(17)(213) <= to_signed(0,32);
  mem_filters(17)(214) <= to_signed(0,32); mem_filters(17)(215) <= to_signed(0,32); mem_filters(17)(216) <= to_signed(0,32);
  mem_filters(17)(217) <= to_signed(0,32); mem_filters(17)(218) <= to_signed(0,32); mem_filters(17)(219) <= to_signed(0,32);
  mem_filters(17)(220) <= to_signed(0,32); mem_filters(17)(221) <= to_signed(0,32); mem_filters(17)(222) <= to_signed(0,32);
  mem_filters(17)(223) <= to_signed(0,32); mem_filters(17)(224) <= to_signed(0,32); mem_filters(17)(225) <= to_signed(0,32);
  mem_filters(17)(226) <= to_signed(0,32); mem_filters(17)(227) <= to_signed(0,32); mem_filters(17)(228) <= to_signed(0,32);
  mem_filters(17)(229) <= to_signed(0,32); mem_filters(17)(230) <= to_signed(0,32); mem_filters(17)(231) <= to_signed(0,32);
  mem_filters(17)(232) <= to_signed(0,32); mem_filters(17)(233) <= to_signed(0,32); mem_filters(17)(234) <= to_signed(0,32);
  mem_filters(17)(235) <= to_signed(0,32); mem_filters(17)(236) <= to_signed(0,32); mem_filters(17)(237) <= to_signed(0,32);
  mem_filters(17)(238) <= to_signed(0,32); mem_filters(17)(239) <= to_signed(0,32); mem_filters(17)(240) <= to_signed(0,32);
  mem_filters(17)(241) <= to_signed(0,32); mem_filters(17)(242) <= to_signed(0,32); mem_filters(17)(243) <= to_signed(0,32);
  mem_filters(17)(244) <= to_signed(0,32); mem_filters(17)(245) <= to_signed(0,32); mem_filters(17)(246) <= to_signed(0,32);
  mem_filters(17)(247) <= to_signed(0,32); mem_filters(17)(248) <= to_signed(0,32); mem_filters(17)(249) <= to_signed(0,32);
  mem_filters(17)(250) <= to_signed(0,32); mem_filters(17)(251) <= to_signed(0,32); mem_filters(17)(252) <= to_signed(0,32);
  mem_filters(17)(253) <= to_signed(0,32); mem_filters(17)(254) <= to_signed(0,32); mem_filters(17)(255) <= to_signed(0,32);
  
  --Filter 18
  mem_filters(18)(0) <= to_signed(0,32); mem_filters(18)(1) <= to_signed(0,32); mem_filters(18)(2) <= to_signed(0,32);
  mem_filters(18)(3) <= to_signed(0,32); mem_filters(18)(4) <= to_signed(0,32); mem_filters(18)(5) <= to_signed(0,32);
  mem_filters(18)(6) <= to_signed(0,32); mem_filters(18)(7) <= to_signed(0,32); mem_filters(18)(8) <= to_signed(0,32);
  mem_filters(18)(9) <= to_signed(0,32); mem_filters(18)(10) <= to_signed(0,32); mem_filters(18)(11) <= to_signed(0,32);
  mem_filters(18)(12) <= to_signed(0,32); mem_filters(18)(13) <= to_signed(0,32); mem_filters(18)(14) <= to_signed(0,32);
  mem_filters(18)(15) <= to_signed(0,32); mem_filters(18)(16) <= to_signed(0,32); mem_filters(18)(17) <= to_signed(0,32);
  mem_filters(18)(18) <= to_signed(0,32); mem_filters(18)(19) <= to_signed(0,32); mem_filters(18)(20) <= to_signed(0,32);
  mem_filters(18)(21) <= to_signed(0,32); mem_filters(18)(22) <= to_signed(0,32); mem_filters(18)(23) <= to_signed(0,32);
  mem_filters(18)(24) <= to_signed(0,32); mem_filters(18)(25) <= to_signed(0,32); mem_filters(18)(26) <= to_signed(0,32);
  mem_filters(18)(27) <= to_signed(0,32); mem_filters(18)(28) <= to_signed(0,32); mem_filters(18)(29) <= to_signed(0,32);
  mem_filters(18)(30) <= to_signed(0,32); mem_filters(18)(31) <= to_signed(0,32); mem_filters(18)(32) <= to_signed(0,32);
  mem_filters(18)(33) <= to_signed(0,32); mem_filters(18)(34) <= to_signed(0,32); mem_filters(18)(35) <= to_signed(0,32);
  mem_filters(18)(36) <= to_signed(0,32); mem_filters(18)(37) <= to_signed(0,32); mem_filters(18)(38) <= to_signed(0,32);
  mem_filters(18)(39) <= to_signed(0,32); mem_filters(18)(40) <= to_signed(0,32); mem_filters(18)(41) <= to_signed(0,32);
  mem_filters(18)(42) <= to_signed(0,32); mem_filters(18)(43) <= to_signed(0,32); mem_filters(18)(44) <= to_signed(0,32);
  mem_filters(18)(45) <= to_signed(0,32);
  mem_filters(18)(46) <= to_signed(0,32); mem_filters(18)(47) <= to_signed(0,32); mem_filters(18)(48) <= to_signed(0,32);
  mem_filters(18)(49) <= to_signed(0,32); mem_filters(18)(50) <= to_signed(0,32); mem_filters(18)(51) <= to_signed(0,32);
  mem_filters(18)(52) <= to_signed(0,32); mem_filters(18)(53) <= to_signed(0,32); mem_filters(18)(54) <= to_signed(0,32);
  mem_filters(18)(55) <= to_signed(0,32); mem_filters(18)(56) <= to_signed(0,32); mem_filters(18)(57) <= to_signed(0,32);
  mem_filters(18)(58) <= to_signed(0,32); mem_filters(18)(59) <= to_signed(0,32); mem_filters(18)(60) <= to_signed(0,32);
  mem_filters(18)(61) <= to_signed(0,32); mem_filters(18)(62) <= to_signed(0,32); mem_filters(18)(63) <= to_signed(0,32);
  mem_filters(18)(64) <= to_signed(0,32); mem_filters(18)(65) <= to_signed(0,32); mem_filters(18)(66) <= to_signed(0,32);
  mem_filters(18)(67) <= to_signed(0,32); mem_filters(18)(68) <= to_signed(0,32); mem_filters(18)(69) <= to_signed(0,32);
  mem_filters(18)(70) <= to_signed(0,32); mem_filters(18)(71) <= to_signed(0,32); mem_filters(18)(72) <= to_signed(0,32);
  mem_filters(18)(73) <= to_signed(0,32); mem_filters(18)(74) <= to_signed(0,32); mem_filters(18)(75) <= to_signed(0,32);
  mem_filters(18)(76) <= to_signed(0,32); mem_filters(18)(77) <= to_signed(0,32); mem_filters(18)(78) <= to_signed(0,32);
  mem_filters(18)(79) <= to_signed(0,32); mem_filters(18)(80) <= to_signed(0,32); mem_filters(18)(81) <= to_signed(0,32);
  mem_filters(18)(82) <= to_signed(0,32); mem_filters(18)(83) <= to_signed(0,32); mem_filters(18)(84) <= to_signed(0,32);
  mem_filters(18)(85) <= to_signed(0,32); mem_filters(18)(86) <= to_signed(0,32); mem_filters(18)(87) <= to_signed(0,32);
  mem_filters(18)(88) <= to_signed(0,32); mem_filters(18)(89) <= to_signed(0,32); mem_filters(18)(90) <= to_signed(0,32);
  mem_filters(18)(91) <= to_signed(0,32); mem_filters(18)(92) <= to_signed(0,32); mem_filters(18)(93) <= to_signed(0,32);
  mem_filters(18)(94) <= to_signed(0,32); mem_filters(18)(95) <= to_signed(0,32); mem_filters(18)(96) <= to_signed(0,32);
  mem_filters(18)(97) <= to_signed(0,32); mem_filters(18)(98) <= to_signed(0,32); mem_filters(18)(99) <= to_signed(0,32);
  mem_filters(18)(100) <= to_signed(0,32); mem_filters(18)(101) <= to_signed(0,32); mem_filters(18)(102) <= to_signed(0,32);
  mem_filters(18)(103) <= to_signed(0,32); mem_filters(18)(104) <= to_signed(0,32); mem_filters(18)(105) <= to_signed(0,32);
  mem_filters(18)(106) <= to_signed(0,32); mem_filters(18)(107) <= to_signed(0,32); mem_filters(18)(108) <= to_signed(0,32);
  mem_filters(18)(109) <= to_signed(0,32); mem_filters(18)(110) <= to_signed(0,32); mem_filters(18)(111) <= to_signed(0,32);
  mem_filters(18)(112) <= to_signed(0,32); mem_filters(18)(113) <= to_signed(0,32); mem_filters(18)(114) <= to_signed(0,32);
  mem_filters(18)(115) <= to_signed(0,32); mem_filters(18)(116) <= to_signed(0,32); mem_filters(18)(117) <= to_signed(0,32);
  mem_filters(18)(118) <= to_signed(0,32); mem_filters(18)(119) <= to_signed(0,32); mem_filters(18)(120) <= to_signed(0,32);
  mem_filters(18)(121) <= to_signed(0,32); mem_filters(18)(122) <= to_signed(0,32); mem_filters(18)(123) <= to_signed(0,32);
  mem_filters(18)(124) <= to_signed(0,32); mem_filters(18)(125) <= to_signed(0,32); mem_filters(18)(126) <= to_signed(0,32);
  mem_filters(18)(127) <= to_signed(0,32); mem_filters(18)(128) <= to_signed(0,32); mem_filters(18)(129) <= to_signed(0,32);
  mem_filters(18)(130) <= to_signed(0,32); mem_filters(18)(131) <= to_signed(0,32); mem_filters(18)(132) <= to_signed(0,32);
  mem_filters(18)(133) <= to_signed(0,32); mem_filters(18)(134) <= to_signed(0,32); mem_filters(18)(135) <= to_signed(0,32);
  mem_filters(18)(136) <= to_signed(0,32); mem_filters(18)(137) <= to_signed(0,32); mem_filters(18)(138) <= to_signed(0,32);
  mem_filters(18)(139) <= to_signed(0,32); mem_filters(18)(140) <= to_signed(0,32); mem_filters(18)(141) <= to_signed(0,32);
  mem_filters(18)(142) <= to_signed(0,32); mem_filters(18)(143) <= to_signed(0,32); mem_filters(18)(144) <= to_signed(0,32);
  mem_filters(18)(145) <= to_signed(0,32); mem_filters(18)(146) <= to_signed(0,32); mem_filters(18)(147) <= to_signed(0,32);
  mem_filters(18)(148) <= to_signed(0,32); mem_filters(18)(149) <= to_signed(0,32); mem_filters(18)(150) <= to_signed(0,32);
  mem_filters(18)(151) <= to_signed(0,32); mem_filters(18)(152) <= to_signed(0,32); mem_filters(18)(153) <= to_signed(0,32);
  mem_filters(18)(154) <= to_signed(0,32); mem_filters(18)(155) <= to_signed(0,32); mem_filters(18)(156) <= to_signed(0,32);
  mem_filters(18)(157) <= to_signed(0,32); mem_filters(18)(158) <= to_signed(0,32); mem_filters(18)(159) <= to_signed(0,32);
  mem_filters(18)(160) <= to_signed(0,32); mem_filters(18)(161) <= to_signed(0,32); mem_filters(18)(162) <= to_signed(0,32);
  mem_filters(18)(163) <= to_signed(0,32); mem_filters(18)(164) <= to_signed(0,32); mem_filters(18)(165) <= to_signed(0,32);
  mem_filters(18)(166) <= to_signed(0,32); mem_filters(18)(167) <= to_signed(0,32); mem_filters(18)(168) <= to_signed(0,32);
  mem_filters(18)(169) <= to_signed(0,32); mem_filters(18)(170) <= to_signed(0,32); mem_filters(18)(171) <= to_signed(0,32);
  mem_filters(18)(172) <= to_signed(0,32); mem_filters(18)(173) <= to_signed(0,32); mem_filters(18)(174) <= to_signed(0,32);
  mem_filters(18)(175) <= to_signed(0,32); mem_filters(18)(176) <= to_signed(0,32); mem_filters(18)(177) <= to_signed(0,32);
  mem_filters(18)(178) <= to_signed(0,32); mem_filters(18)(179) <= to_signed(0,32); mem_filters(18)(180) <= to_signed(0,32);
  mem_filters(18)(181) <= to_signed(0,32); mem_filters(18)(182) <= to_signed(0,32); mem_filters(18)(183) <= to_signed(0,32);
  mem_filters(18)(184) <= to_signed(0,32); mem_filters(18)(185) <= to_signed(0,32); mem_filters(18)(186) <= to_signed(0,32);
  mem_filters(18)(187) <= to_signed(0,32); mem_filters(18)(188) <= to_signed(0,32); mem_filters(18)(189) <= to_signed(0,32);
  mem_filters(18)(190) <= to_signed(0,32); mem_filters(18)(191) <= to_signed(0,32); mem_filters(18)(192) <= to_signed(0,32);
  mem_filters(18)(193) <= to_signed(0,32); mem_filters(18)(194) <= to_signed(0,32); mem_filters(18)(195) <= to_signed(0,32);
  mem_filters(18)(196) <= to_signed(0,32); mem_filters(18)(197) <= to_signed(0,32); mem_filters(18)(198) <= to_signed(0,32);
  mem_filters(18)(199) <= to_signed(0,32); mem_filters(18)(200) <= to_signed(0,32); mem_filters(18)(201) <= to_signed(0,32);
  mem_filters(18)(202) <= to_signed(0,32); mem_filters(18)(203) <= to_signed(0,32); mem_filters(18)(204) <= to_signed(0,32);
  mem_filters(18)(205) <= to_signed(0,32); mem_filters(18)(206) <= to_signed(0,32); mem_filters(18)(207) <= to_signed(0,32);
  mem_filters(18)(208) <= to_signed(0,32); mem_filters(18)(209) <= to_signed(0,32); mem_filters(18)(210) <= to_signed(0,32);
  mem_filters(18)(211) <= to_signed(0,32); mem_filters(18)(212) <= to_signed(0,32); mem_filters(18)(213) <= to_signed(0,32);
  mem_filters(18)(214) <= to_signed(0,32); mem_filters(18)(215) <= to_signed(0,32); mem_filters(18)(216) <= to_signed(0,32);
  mem_filters(18)(217) <= to_signed(0,32); mem_filters(18)(218) <= to_signed(0,32); mem_filters(18)(219) <= to_signed(0,32);
  mem_filters(18)(220) <= to_signed(0,32); mem_filters(18)(221) <= to_signed(0,32); mem_filters(18)(222) <= to_signed(0,32);
  mem_filters(18)(223) <= to_signed(0,32); mem_filters(18)(224) <= to_signed(0,32); mem_filters(18)(225) <= to_signed(0,32);
  mem_filters(18)(226) <= to_signed(0,32); mem_filters(18)(227) <= to_signed(0,32); mem_filters(18)(228) <= to_signed(0,32);
  mem_filters(18)(229) <= to_signed(0,32); mem_filters(18)(230) <= to_signed(0,32); mem_filters(18)(231) <= to_signed(0,32);
  mem_filters(18)(232) <= to_signed(0,32); mem_filters(18)(233) <= to_signed(0,32); mem_filters(18)(234) <= to_signed(0,32);
  mem_filters(18)(235) <= to_signed(0,32); mem_filters(18)(236) <= to_signed(0,32); mem_filters(18)(237) <= to_signed(0,32);
  mem_filters(18)(238) <= to_signed(0,32); mem_filters(18)(239) <= to_signed(0,32); mem_filters(18)(240) <= to_signed(0,32);
  mem_filters(18)(241) <= to_signed(0,32); mem_filters(18)(242) <= to_signed(0,32); mem_filters(18)(243) <= to_signed(0,32);
  mem_filters(18)(244) <= to_signed(0,32); mem_filters(18)(245) <= to_signed(0,32); mem_filters(18)(246) <= to_signed(0,32);
  mem_filters(18)(247) <= to_signed(0,32); mem_filters(18)(248) <= to_signed(0,32); mem_filters(18)(249) <= to_signed(0,32);
  mem_filters(18)(250) <= to_signed(0,32); mem_filters(18)(251) <= to_signed(0,32); mem_filters(18)(252) <= to_signed(0,32);
  mem_filters(18)(253) <= to_signed(0,32); mem_filters(18)(254) <= to_signed(0,32); mem_filters(18)(255) <= to_signed(0,32);
  
  --Filter 19
  mem_filters(19)(0) <= to_signed(0,32); mem_filters(19)(1) <= to_signed(0,32); mem_filters(19)(2) <= to_signed(0,32);
  mem_filters(19)(3) <= to_signed(0,32); mem_filters(19)(4) <= to_signed(0,32); mem_filters(19)(5) <= to_signed(0,32);
  mem_filters(19)(6) <= to_signed(0,32); mem_filters(19)(7) <= to_signed(0,32); mem_filters(19)(8) <= to_signed(0,32);
  mem_filters(19)(9) <= to_signed(0,32); mem_filters(19)(10) <= to_signed(0,32); mem_filters(19)(11) <= to_signed(0,32);
  mem_filters(19)(12) <= to_signed(0,32); mem_filters(19)(13) <= to_signed(0,32); mem_filters(19)(14) <= to_signed(0,32);
  mem_filters(19)(15) <= to_signed(0,32); mem_filters(19)(16) <= to_signed(0,32); mem_filters(19)(17) <= to_signed(0,32);
  mem_filters(19)(18) <= to_signed(0,32); mem_filters(19)(19) <= to_signed(0,32); mem_filters(19)(20) <= to_signed(0,32);
  mem_filters(19)(21) <= to_signed(0,32); mem_filters(19)(22) <= to_signed(0,32); mem_filters(19)(23) <= to_signed(0,32);
  mem_filters(19)(24) <= to_signed(0,32); mem_filters(19)(25) <= to_signed(0,32); mem_filters(19)(26) <= to_signed(0,32);
  mem_filters(19)(27) <= to_signed(0,32); mem_filters(19)(28) <= to_signed(0,32); mem_filters(19)(29) <= to_signed(0,32);
  mem_filters(19)(30) <= to_signed(0,32); mem_filters(19)(31) <= to_signed(0,32); mem_filters(19)(32) <= to_signed(0,32);
  mem_filters(19)(33) <= to_signed(0,32); mem_filters(19)(34) <= to_signed(0,32); mem_filters(19)(35) <= to_signed(0,32);
  mem_filters(19)(36) <= to_signed(0,32); mem_filters(19)(37) <= to_signed(0,32); mem_filters(19)(38) <= to_signed(0,32);
  mem_filters(19)(39) <= to_signed(0,32); mem_filters(19)(40) <= to_signed(0,32); mem_filters(19)(41) <= to_signed(0,32);
  mem_filters(19)(42) <= to_signed(0,32); mem_filters(19)(43) <= to_signed(0,32); mem_filters(19)(44) <= to_signed(0,32);
  mem_filters(19)(45) <= to_signed(0,32);
  mem_filters(19)(46) <= to_signed(0,32); mem_filters(19)(47) <= to_signed(0,32); mem_filters(19)(48) <= to_signed(0,32);
  mem_filters(19)(49) <= to_signed(0,32); mem_filters(19)(50) <= to_signed(0,32); mem_filters(19)(51) <= to_signed(0,32);
  mem_filters(19)(52) <= to_signed(0,32); mem_filters(19)(53) <= to_signed(0,32); mem_filters(19)(54) <= to_signed(0,32);
  mem_filters(19)(55) <= to_signed(0,32); mem_filters(19)(56) <= to_signed(0,32); mem_filters(19)(57) <= to_signed(0,32);
  mem_filters(19)(58) <= to_signed(0,32); mem_filters(19)(59) <= to_signed(0,32); mem_filters(19)(60) <= to_signed(0,32);
  mem_filters(19)(61) <= to_signed(0,32); mem_filters(19)(62) <= to_signed(0,32); mem_filters(19)(63) <= to_signed(0,32);
  mem_filters(19)(64) <= to_signed(0,32); mem_filters(19)(65) <= to_signed(0,32); mem_filters(19)(66) <= to_signed(0,32);
  mem_filters(19)(67) <= to_signed(0,32); mem_filters(19)(68) <= to_signed(0,32); mem_filters(19)(69) <= to_signed(0,32);
  mem_filters(19)(70) <= to_signed(0,32); mem_filters(19)(71) <= to_signed(0,32); mem_filters(19)(72) <= to_signed(0,32);
  mem_filters(19)(73) <= to_signed(0,32); mem_filters(19)(74) <= to_signed(0,32); mem_filters(19)(75) <= to_signed(0,32);
  mem_filters(19)(76) <= to_signed(0,32); mem_filters(19)(77) <= to_signed(0,32); mem_filters(19)(78) <= to_signed(0,32);
  mem_filters(19)(79) <= to_signed(0,32); mem_filters(19)(80) <= to_signed(0,32); mem_filters(19)(81) <= to_signed(0,32);
  mem_filters(19)(82) <= to_signed(0,32); mem_filters(19)(83) <= to_signed(0,32); mem_filters(19)(84) <= to_signed(0,32);
  mem_filters(19)(85) <= to_signed(0,32); mem_filters(19)(86) <= to_signed(0,32); mem_filters(19)(87) <= to_signed(0,32);
  mem_filters(19)(88) <= to_signed(0,32); mem_filters(19)(89) <= to_signed(0,32); mem_filters(19)(90) <= to_signed(0,32);
  mem_filters(19)(91) <= to_signed(0,32); mem_filters(19)(92) <= to_signed(0,32); mem_filters(19)(93) <= to_signed(0,32);
  mem_filters(19)(94) <= to_signed(0,32); mem_filters(19)(95) <= to_signed(0,32); mem_filters(19)(96) <= to_signed(0,32);
  mem_filters(19)(97) <= to_signed(0,32); mem_filters(19)(98) <= to_signed(0,32); mem_filters(19)(99) <= to_signed(0,32);
  mem_filters(19)(100) <= to_signed(0,32); mem_filters(19)(101) <= to_signed(0,32); mem_filters(19)(102) <= to_signed(0,32);
  mem_filters(19)(103) <= to_signed(0,32); mem_filters(19)(104) <= to_signed(0,32); mem_filters(19)(105) <= to_signed(0,32);
  mem_filters(19)(106) <= to_signed(0,32); mem_filters(19)(107) <= to_signed(0,32); mem_filters(19)(108) <= to_signed(0,32);
  mem_filters(19)(109) <= to_signed(0,32); mem_filters(19)(110) <= to_signed(0,32); mem_filters(19)(111) <= to_signed(0,32);
  mem_filters(19)(112) <= to_signed(0,32); mem_filters(19)(113) <= to_signed(0,32); mem_filters(19)(114) <= to_signed(0,32);
  mem_filters(19)(115) <= to_signed(0,32); mem_filters(19)(116) <= to_signed(0,32); mem_filters(19)(117) <= to_signed(0,32);
  mem_filters(19)(118) <= to_signed(0,32); mem_filters(19)(119) <= to_signed(0,32); mem_filters(19)(120) <= to_signed(0,32);
  mem_filters(19)(121) <= to_signed(0,32); mem_filters(19)(122) <= to_signed(0,32); mem_filters(19)(123) <= to_signed(0,32);
  mem_filters(19)(124) <= to_signed(0,32); mem_filters(19)(125) <= to_signed(0,32); mem_filters(19)(126) <= to_signed(0,32);
  mem_filters(19)(127) <= to_signed(0,32); mem_filters(19)(128) <= to_signed(0,32); mem_filters(19)(129) <= to_signed(0,32);
  mem_filters(19)(130) <= to_signed(0,32); mem_filters(19)(131) <= to_signed(0,32); mem_filters(19)(132) <= to_signed(0,32);
  mem_filters(19)(133) <= to_signed(0,32); mem_filters(19)(134) <= to_signed(0,32); mem_filters(19)(135) <= to_signed(0,32);
  mem_filters(19)(136) <= to_signed(0,32); mem_filters(19)(137) <= to_signed(0,32); mem_filters(19)(138) <= to_signed(0,32);
  mem_filters(19)(139) <= to_signed(0,32); mem_filters(19)(140) <= to_signed(0,32); mem_filters(19)(141) <= to_signed(0,32);
  mem_filters(19)(142) <= to_signed(0,32); mem_filters(19)(143) <= to_signed(0,32); mem_filters(19)(144) <= to_signed(0,32);
  mem_filters(19)(145) <= to_signed(0,32); mem_filters(19)(146) <= to_signed(0,32); mem_filters(19)(147) <= to_signed(0,32);
  mem_filters(19)(148) <= to_signed(0,32); mem_filters(19)(149) <= to_signed(0,32); mem_filters(19)(150) <= to_signed(0,32);
  mem_filters(19)(151) <= to_signed(0,32); mem_filters(19)(152) <= to_signed(0,32); mem_filters(19)(153) <= to_signed(0,32);
  mem_filters(19)(154) <= to_signed(0,32); mem_filters(19)(155) <= to_signed(0,32); mem_filters(19)(156) <= to_signed(0,32);
  mem_filters(19)(157) <= to_signed(0,32); mem_filters(19)(158) <= to_signed(0,32); mem_filters(19)(159) <= to_signed(0,32);
  mem_filters(19)(160) <= to_signed(0,32); mem_filters(19)(161) <= to_signed(0,32); mem_filters(19)(162) <= to_signed(0,32);
  mem_filters(19)(163) <= to_signed(0,32); mem_filters(19)(164) <= to_signed(0,32); mem_filters(19)(165) <= to_signed(0,32);
  mem_filters(19)(166) <= to_signed(0,32); mem_filters(19)(167) <= to_signed(0,32); mem_filters(19)(168) <= to_signed(0,32);
  mem_filters(19)(169) <= to_signed(0,32); mem_filters(19)(170) <= to_signed(0,32); mem_filters(19)(171) <= to_signed(0,32);
  mem_filters(19)(172) <= to_signed(0,32); mem_filters(19)(173) <= to_signed(0,32); mem_filters(19)(174) <= to_signed(0,32);
  mem_filters(19)(175) <= to_signed(0,32); mem_filters(19)(176) <= to_signed(0,32); mem_filters(19)(177) <= to_signed(0,32);
  mem_filters(19)(178) <= to_signed(0,32); mem_filters(19)(179) <= to_signed(0,32); mem_filters(19)(180) <= to_signed(0,32);
  mem_filters(19)(181) <= to_signed(0,32); mem_filters(19)(182) <= to_signed(0,32); mem_filters(19)(183) <= to_signed(0,32);
  mem_filters(19)(184) <= to_signed(0,32); mem_filters(19)(185) <= to_signed(0,32); mem_filters(19)(186) <= to_signed(0,32);
  mem_filters(19)(187) <= to_signed(0,32); mem_filters(19)(188) <= to_signed(0,32); mem_filters(19)(189) <= to_signed(0,32);
  mem_filters(19)(190) <= to_signed(0,32); mem_filters(19)(191) <= to_signed(0,32); mem_filters(19)(192) <= to_signed(0,32);
  mem_filters(19)(193) <= to_signed(0,32); mem_filters(19)(194) <= to_signed(0,32); mem_filters(19)(195) <= to_signed(0,32);
  mem_filters(19)(196) <= to_signed(0,32); mem_filters(19)(197) <= to_signed(0,32); mem_filters(19)(198) <= to_signed(0,32);
  mem_filters(19)(199) <= to_signed(0,32); mem_filters(19)(200) <= to_signed(0,32); mem_filters(19)(201) <= to_signed(0,32);
  mem_filters(19)(202) <= to_signed(0,32); mem_filters(19)(203) <= to_signed(0,32); mem_filters(19)(204) <= to_signed(0,32);
  mem_filters(19)(205) <= to_signed(0,32); mem_filters(19)(206) <= to_signed(0,32); mem_filters(19)(207) <= to_signed(0,32);
  mem_filters(19)(208) <= to_signed(0,32); mem_filters(19)(209) <= to_signed(0,32); mem_filters(19)(210) <= to_signed(0,32);
  mem_filters(19)(211) <= to_signed(0,32); mem_filters(19)(212) <= to_signed(0,32); mem_filters(19)(213) <= to_signed(0,32);
  mem_filters(19)(214) <= to_signed(0,32); mem_filters(19)(215) <= to_signed(0,32); mem_filters(19)(216) <= to_signed(0,32);
  mem_filters(19)(217) <= to_signed(0,32); mem_filters(19)(218) <= to_signed(0,32); mem_filters(19)(219) <= to_signed(0,32);
  mem_filters(19)(220) <= to_signed(0,32); mem_filters(19)(221) <= to_signed(0,32); mem_filters(19)(222) <= to_signed(0,32);
  mem_filters(19)(223) <= to_signed(0,32); mem_filters(19)(224) <= to_signed(0,32); mem_filters(19)(225) <= to_signed(0,32);
  mem_filters(19)(226) <= to_signed(0,32); mem_filters(19)(227) <= to_signed(0,32); mem_filters(19)(228) <= to_signed(0,32);
  mem_filters(19)(229) <= to_signed(0,32); mem_filters(19)(230) <= to_signed(0,32); mem_filters(19)(231) <= to_signed(0,32);
  mem_filters(19)(232) <= to_signed(0,32); mem_filters(19)(233) <= to_signed(0,32); mem_filters(19)(234) <= to_signed(0,32);
  mem_filters(19)(235) <= to_signed(0,32); mem_filters(19)(236) <= to_signed(0,32); mem_filters(19)(237) <= to_signed(0,32);
  mem_filters(19)(238) <= to_signed(0,32); mem_filters(19)(239) <= to_signed(0,32); mem_filters(19)(240) <= to_signed(0,32);
  mem_filters(19)(241) <= to_signed(0,32); mem_filters(19)(242) <= to_signed(0,32); mem_filters(19)(243) <= to_signed(0,32);
  mem_filters(19)(244) <= to_signed(0,32); mem_filters(19)(245) <= to_signed(0,32); mem_filters(19)(246) <= to_signed(0,32);
  mem_filters(19)(247) <= to_signed(0,32); mem_filters(19)(248) <= to_signed(0,32); mem_filters(19)(249) <= to_signed(0,32);
  mem_filters(19)(250) <= to_signed(0,32); mem_filters(19)(251) <= to_signed(0,32); mem_filters(19)(252) <= to_signed(0,32);
  mem_filters(19)(253) <= to_signed(0,32); mem_filters(19)(254) <= to_signed(0,32); mem_filters(19)(255) <= to_signed(0,32);
  
  --Filter 20
  mem_filters(20)(0) <= to_signed(0,32); mem_filters(20)(1) <= to_signed(0,32); mem_filters(20)(2) <= to_signed(0,32);
  mem_filters(20)(3) <= to_signed(0,32); mem_filters(20)(4) <= to_signed(0,32); mem_filters(20)(5) <= to_signed(0,32);
  mem_filters(20)(6) <= to_signed(0,32); mem_filters(20)(7) <= to_signed(0,32); mem_filters(20)(8) <= to_signed(0,32);
  mem_filters(20)(9) <= to_signed(0,32); mem_filters(20)(10) <= to_signed(0,32); mem_filters(20)(11) <= to_signed(0,32);
  mem_filters(20)(12) <= to_signed(0,32); mem_filters(20)(13) <= to_signed(0,32); mem_filters(20)(14) <= to_signed(0,32);
  mem_filters(20)(15) <= to_signed(0,32); mem_filters(20)(16) <= to_signed(0,32); mem_filters(20)(17) <= to_signed(0,32);
  mem_filters(20)(18) <= to_signed(0,32); mem_filters(20)(19) <= to_signed(0,32); mem_filters(20)(20) <= to_signed(0,32);
  mem_filters(20)(21) <= to_signed(0,32); mem_filters(20)(22) <= to_signed(0,32); mem_filters(20)(23) <= to_signed(0,32);
  mem_filters(20)(24) <= to_signed(0,32); mem_filters(20)(25) <= to_signed(0,32); mem_filters(20)(26) <= to_signed(0,32);
  mem_filters(20)(27) <= to_signed(0,32); mem_filters(20)(28) <= to_signed(0,32); mem_filters(20)(29) <= to_signed(0,32);
  mem_filters(20)(30) <= to_signed(0,32); mem_filters(20)(31) <= to_signed(0,32); mem_filters(20)(32) <= to_signed(0,32);
  mem_filters(20)(33) <= to_signed(0,32); mem_filters(20)(34) <= to_signed(0,32); mem_filters(20)(35) <= to_signed(0,32);
  mem_filters(20)(36) <= to_signed(0,32); mem_filters(20)(37) <= to_signed(0,32); mem_filters(20)(38) <= to_signed(0,32);
  mem_filters(20)(39) <= to_signed(0,32); mem_filters(20)(40) <= to_signed(0,32); mem_filters(20)(41) <= to_signed(0,32);
  mem_filters(20)(42) <= to_signed(0,32); mem_filters(20)(43) <= to_signed(0,32); mem_filters(20)(44) <= to_signed(0,32);
  mem_filters(20)(45) <= to_signed(0,32);
  mem_filters(20)(46) <= to_signed(0,32); mem_filters(20)(47) <= to_signed(0,32); mem_filters(20)(48) <= to_signed(0,32);
  mem_filters(20)(49) <= to_signed(0,32); mem_filters(20)(50) <= to_signed(0,32); mem_filters(20)(51) <= to_signed(0,32);
  mem_filters(20)(52) <= to_signed(0,32); mem_filters(20)(53) <= to_signed(0,32); mem_filters(20)(54) <= to_signed(0,32);
  mem_filters(20)(55) <= to_signed(0,32); mem_filters(20)(56) <= to_signed(0,32); mem_filters(20)(57) <= to_signed(0,32);
  mem_filters(20)(58) <= to_signed(0,32); mem_filters(20)(59) <= to_signed(0,32); mem_filters(20)(60) <= to_signed(0,32);
  mem_filters(20)(61) <= to_signed(0,32); mem_filters(20)(62) <= to_signed(0,32); mem_filters(20)(63) <= to_signed(0,32);
  mem_filters(20)(64) <= to_signed(0,32); mem_filters(20)(65) <= to_signed(0,32); mem_filters(20)(66) <= to_signed(0,32);
  mem_filters(20)(67) <= to_signed(0,32); mem_filters(20)(68) <= to_signed(0,32); mem_filters(20)(69) <= to_signed(0,32);
  mem_filters(20)(70) <= to_signed(0,32); mem_filters(20)(71) <= to_signed(0,32); mem_filters(20)(72) <= to_signed(0,32);
  mem_filters(20)(73) <= to_signed(0,32); mem_filters(20)(74) <= to_signed(0,32); mem_filters(20)(75) <= to_signed(0,32);
  mem_filters(20)(76) <= to_signed(0,32); mem_filters(20)(77) <= to_signed(0,32); mem_filters(20)(78) <= to_signed(0,32);
  mem_filters(20)(79) <= to_signed(0,32); mem_filters(20)(80) <= to_signed(0,32); mem_filters(20)(81) <= to_signed(0,32);
  mem_filters(20)(82) <= to_signed(0,32); mem_filters(20)(83) <= to_signed(0,32); mem_filters(20)(84) <= to_signed(0,32);
  mem_filters(20)(85) <= to_signed(0,32); mem_filters(20)(86) <= to_signed(0,32); mem_filters(20)(87) <= to_signed(0,32);
  mem_filters(20)(88) <= to_signed(0,32); mem_filters(20)(89) <= to_signed(0,32); mem_filters(20)(90) <= to_signed(0,32);
  mem_filters(20)(91) <= to_signed(0,32); mem_filters(20)(92) <= to_signed(0,32); mem_filters(20)(93) <= to_signed(0,32);
  mem_filters(20)(94) <= to_signed(0,32); mem_filters(20)(95) <= to_signed(0,32); mem_filters(20)(96) <= to_signed(0,32);
  mem_filters(20)(97) <= to_signed(0,32); mem_filters(20)(98) <= to_signed(0,32); mem_filters(20)(99) <= to_signed(0,32);
  mem_filters(20)(100) <= to_signed(0,32); mem_filters(20)(101) <= to_signed(0,32); mem_filters(20)(102) <= to_signed(0,32);
  mem_filters(20)(103) <= to_signed(0,32); mem_filters(20)(104) <= to_signed(0,32); mem_filters(20)(105) <= to_signed(0,32);
  mem_filters(20)(106) <= to_signed(0,32); mem_filters(20)(107) <= to_signed(0,32); mem_filters(20)(108) <= to_signed(0,32);
  mem_filters(20)(109) <= to_signed(0,32); mem_filters(20)(110) <= to_signed(0,32); mem_filters(20)(111) <= to_signed(0,32);
  mem_filters(20)(112) <= to_signed(0,32); mem_filters(20)(113) <= to_signed(0,32); mem_filters(20)(114) <= to_signed(0,32);
  mem_filters(20)(115) <= to_signed(0,32); mem_filters(20)(116) <= to_signed(0,32); mem_filters(20)(117) <= to_signed(0,32);
  mem_filters(20)(118) <= to_signed(0,32); mem_filters(20)(119) <= to_signed(0,32); mem_filters(20)(120) <= to_signed(0,32);
  mem_filters(20)(121) <= to_signed(0,32); mem_filters(20)(122) <= to_signed(0,32); mem_filters(20)(123) <= to_signed(0,32);
  mem_filters(20)(124) <= to_signed(0,32); mem_filters(20)(125) <= to_signed(0,32); mem_filters(20)(126) <= to_signed(0,32);
  mem_filters(20)(127) <= to_signed(0,32); mem_filters(20)(128) <= to_signed(0,32); mem_filters(20)(129) <= to_signed(0,32);
  mem_filters(20)(130) <= to_signed(0,32); mem_filters(20)(131) <= to_signed(0,32); mem_filters(20)(132) <= to_signed(0,32);
  mem_filters(20)(133) <= to_signed(0,32); mem_filters(20)(134) <= to_signed(0,32); mem_filters(20)(135) <= to_signed(0,32);
  mem_filters(20)(136) <= to_signed(0,32); mem_filters(20)(137) <= to_signed(0,32); mem_filters(20)(138) <= to_signed(0,32);
  mem_filters(20)(139) <= to_signed(0,32); mem_filters(20)(140) <= to_signed(0,32); mem_filters(20)(141) <= to_signed(0,32);
  mem_filters(20)(142) <= to_signed(0,32); mem_filters(20)(143) <= to_signed(0,32); mem_filters(20)(144) <= to_signed(0,32);
  mem_filters(20)(145) <= to_signed(0,32); mem_filters(20)(146) <= to_signed(0,32); mem_filters(20)(147) <= to_signed(0,32);
  mem_filters(20)(148) <= to_signed(0,32); mem_filters(20)(149) <= to_signed(0,32); mem_filters(20)(150) <= to_signed(0,32);
  mem_filters(20)(151) <= to_signed(0,32); mem_filters(20)(152) <= to_signed(0,32); mem_filters(20)(153) <= to_signed(0,32);
  mem_filters(20)(154) <= to_signed(0,32); mem_filters(20)(155) <= to_signed(0,32); mem_filters(20)(156) <= to_signed(0,32);
  mem_filters(20)(157) <= to_signed(0,32); mem_filters(20)(158) <= to_signed(0,32); mem_filters(20)(159) <= to_signed(0,32);
  mem_filters(20)(160) <= to_signed(0,32); mem_filters(20)(161) <= to_signed(0,32); mem_filters(20)(162) <= to_signed(0,32);
  mem_filters(20)(163) <= to_signed(0,32); mem_filters(20)(164) <= to_signed(0,32); mem_filters(20)(165) <= to_signed(0,32);
  mem_filters(20)(166) <= to_signed(0,32); mem_filters(20)(167) <= to_signed(0,32); mem_filters(20)(168) <= to_signed(0,32);
  mem_filters(20)(169) <= to_signed(0,32); mem_filters(20)(170) <= to_signed(0,32); mem_filters(20)(171) <= to_signed(0,32);
  mem_filters(20)(172) <= to_signed(0,32); mem_filters(20)(173) <= to_signed(0,32); mem_filters(20)(174) <= to_signed(0,32);
  mem_filters(20)(175) <= to_signed(0,32); mem_filters(20)(176) <= to_signed(0,32); mem_filters(20)(177) <= to_signed(0,32);
  mem_filters(20)(178) <= to_signed(0,32); mem_filters(20)(179) <= to_signed(0,32); mem_filters(20)(180) <= to_signed(0,32);
  mem_filters(20)(181) <= to_signed(0,32); mem_filters(20)(182) <= to_signed(0,32); mem_filters(20)(183) <= to_signed(0,32);
  mem_filters(20)(184) <= to_signed(0,32); mem_filters(20)(185) <= to_signed(0,32); mem_filters(20)(186) <= to_signed(0,32);
  mem_filters(20)(187) <= to_signed(0,32); mem_filters(20)(188) <= to_signed(0,32); mem_filters(20)(189) <= to_signed(0,32);
  mem_filters(20)(190) <= to_signed(0,32); mem_filters(20)(191) <= to_signed(0,32); mem_filters(20)(192) <= to_signed(0,32);
  mem_filters(20)(193) <= to_signed(0,32); mem_filters(20)(194) <= to_signed(0,32); mem_filters(20)(195) <= to_signed(0,32);
  mem_filters(20)(196) <= to_signed(0,32); mem_filters(20)(197) <= to_signed(0,32); mem_filters(20)(198) <= to_signed(0,32);
  mem_filters(20)(199) <= to_signed(0,32); mem_filters(20)(200) <= to_signed(0,32); mem_filters(20)(201) <= to_signed(0,32);
  mem_filters(20)(202) <= to_signed(0,32); mem_filters(20)(203) <= to_signed(0,32); mem_filters(20)(204) <= to_signed(0,32);
  mem_filters(20)(205) <= to_signed(0,32); mem_filters(20)(206) <= to_signed(0,32); mem_filters(20)(207) <= to_signed(0,32);
  mem_filters(20)(208) <= to_signed(0,32); mem_filters(20)(209) <= to_signed(0,32); mem_filters(20)(210) <= to_signed(0,32);
  mem_filters(20)(211) <= to_signed(0,32); mem_filters(20)(212) <= to_signed(0,32); mem_filters(20)(213) <= to_signed(0,32);
  mem_filters(20)(214) <= to_signed(0,32); mem_filters(20)(215) <= to_signed(0,32); mem_filters(20)(216) <= to_signed(0,32);
  mem_filters(20)(217) <= to_signed(0,32); mem_filters(20)(218) <= to_signed(0,32); mem_filters(20)(219) <= to_signed(0,32);
  mem_filters(20)(220) <= to_signed(0,32); mem_filters(20)(221) <= to_signed(0,32); mem_filters(20)(222) <= to_signed(0,32);
  mem_filters(20)(223) <= to_signed(0,32); mem_filters(20)(224) <= to_signed(0,32); mem_filters(20)(225) <= to_signed(0,32);
  mem_filters(20)(226) <= to_signed(0,32); mem_filters(20)(227) <= to_signed(0,32); mem_filters(20)(228) <= to_signed(0,32);
  mem_filters(20)(229) <= to_signed(0,32); mem_filters(20)(230) <= to_signed(0,32); mem_filters(20)(231) <= to_signed(0,32);
  mem_filters(20)(232) <= to_signed(0,32); mem_filters(20)(233) <= to_signed(0,32); mem_filters(20)(234) <= to_signed(0,32);
  mem_filters(20)(235) <= to_signed(0,32); mem_filters(20)(236) <= to_signed(0,32); mem_filters(20)(237) <= to_signed(0,32);
  mem_filters(20)(238) <= to_signed(0,32); mem_filters(20)(239) <= to_signed(0,32); mem_filters(20)(240) <= to_signed(0,32);
  mem_filters(20)(241) <= to_signed(0,32); mem_filters(20)(242) <= to_signed(0,32); mem_filters(20)(243) <= to_signed(0,32);
  mem_filters(20)(244) <= to_signed(0,32); mem_filters(20)(245) <= to_signed(0,32); mem_filters(20)(246) <= to_signed(0,32);
  mem_filters(20)(247) <= to_signed(0,32); mem_filters(20)(248) <= to_signed(0,32); mem_filters(20)(249) <= to_signed(0,32);
  mem_filters(20)(250) <= to_signed(0,32); mem_filters(20)(251) <= to_signed(0,32); mem_filters(20)(252) <= to_signed(0,32);
  mem_filters(20)(253) <= to_signed(0,32); mem_filters(20)(254) <= to_signed(0,32); mem_filters(20)(255) <= to_signed(0,32);
  
  --Filter 21
  mem_filters(21)(0) <= to_signed(0,32); mem_filters(21)(1) <= to_signed(0,32); mem_filters(21)(2) <= to_signed(0,32);
  mem_filters(21)(3) <= to_signed(0,32); mem_filters(21)(4) <= to_signed(0,32); mem_filters(21)(5) <= to_signed(0,32);
  mem_filters(21)(6) <= to_signed(0,32); mem_filters(21)(7) <= to_signed(0,32); mem_filters(21)(8) <= to_signed(0,32);
  mem_filters(21)(9) <= to_signed(0,32); mem_filters(21)(10) <= to_signed(0,32); mem_filters(21)(11) <= to_signed(0,32);
  mem_filters(21)(12) <= to_signed(0,32); mem_filters(21)(13) <= to_signed(0,32); mem_filters(21)(14) <= to_signed(0,32);
  mem_filters(21)(15) <= to_signed(0,32); mem_filters(21)(16) <= to_signed(0,32); mem_filters(21)(17) <= to_signed(0,32);
  mem_filters(21)(18) <= to_signed(0,32); mem_filters(21)(19) <= to_signed(0,32); mem_filters(21)(20) <= to_signed(0,32);
  mem_filters(21)(21) <= to_signed(0,32); mem_filters(21)(22) <= to_signed(0,32); mem_filters(21)(23) <= to_signed(0,32);
  mem_filters(21)(24) <= to_signed(0,32); mem_filters(21)(25) <= to_signed(0,32); mem_filters(21)(26) <= to_signed(0,32);
  mem_filters(21)(27) <= to_signed(0,32); mem_filters(21)(28) <= to_signed(0,32); mem_filters(21)(29) <= to_signed(0,32);
  mem_filters(21)(30) <= to_signed(0,32); mem_filters(21)(31) <= to_signed(0,32); mem_filters(21)(32) <= to_signed(0,32);
  mem_filters(21)(33) <= to_signed(0,32); mem_filters(21)(34) <= to_signed(0,32); mem_filters(21)(35) <= to_signed(0,32);
  mem_filters(21)(36) <= to_signed(0,32); mem_filters(21)(37) <= to_signed(0,32); mem_filters(21)(38) <= to_signed(0,32);
  mem_filters(21)(39) <= to_signed(0,32); mem_filters(21)(40) <= to_signed(0,32); mem_filters(21)(41) <= to_signed(0,32);
  mem_filters(21)(42) <= to_signed(0,32); mem_filters(21)(43) <= to_signed(0,32); mem_filters(21)(44) <= to_signed(0,32);
  mem_filters(21)(45) <= to_signed(0,32);
  mem_filters(21)(46) <= to_signed(0,32); mem_filters(21)(47) <= to_signed(0,32); mem_filters(21)(48) <= to_signed(0,32);
  mem_filters(21)(49) <= to_signed(0,32); mem_filters(21)(50) <= to_signed(0,32); mem_filters(21)(51) <= to_signed(0,32);
  mem_filters(21)(52) <= to_signed(0,32); mem_filters(21)(53) <= to_signed(0,32); mem_filters(21)(54) <= to_signed(0,32);
  mem_filters(21)(55) <= to_signed(0,32); mem_filters(21)(56) <= to_signed(0,32); mem_filters(21)(57) <= to_signed(0,32);
  mem_filters(21)(58) <= to_signed(0,32); mem_filters(21)(59) <= to_signed(0,32); mem_filters(21)(60) <= to_signed(0,32);
  mem_filters(21)(61) <= to_signed(0,32); mem_filters(21)(62) <= to_signed(0,32); mem_filters(21)(63) <= to_signed(0,32);
  mem_filters(21)(64) <= to_signed(0,32); mem_filters(21)(65) <= to_signed(0,32); mem_filters(21)(66) <= to_signed(0,32);
  mem_filters(21)(67) <= to_signed(0,32); mem_filters(21)(68) <= to_signed(0,32); mem_filters(21)(69) <= to_signed(0,32);
  mem_filters(21)(70) <= to_signed(0,32); mem_filters(21)(71) <= to_signed(0,32); mem_filters(21)(72) <= to_signed(0,32);
  mem_filters(21)(73) <= to_signed(0,32); mem_filters(21)(74) <= to_signed(0,32); mem_filters(21)(75) <= to_signed(0,32);
  mem_filters(21)(76) <= to_signed(0,32); mem_filters(21)(77) <= to_signed(0,32); mem_filters(21)(78) <= to_signed(0,32);
  mem_filters(21)(79) <= to_signed(0,32); mem_filters(21)(80) <= to_signed(0,32); mem_filters(21)(81) <= to_signed(0,32);
  mem_filters(21)(82) <= to_signed(0,32); mem_filters(21)(83) <= to_signed(0,32); mem_filters(21)(84) <= to_signed(0,32);
  mem_filters(21)(85) <= to_signed(0,32); mem_filters(21)(86) <= to_signed(0,32); mem_filters(21)(87) <= to_signed(0,32);
  mem_filters(21)(88) <= to_signed(0,32); mem_filters(21)(89) <= to_signed(0,32); mem_filters(21)(90) <= to_signed(0,32);
  mem_filters(21)(91) <= to_signed(0,32); mem_filters(21)(92) <= to_signed(0,32); mem_filters(21)(93) <= to_signed(0,32);
  mem_filters(21)(94) <= to_signed(0,32); mem_filters(21)(95) <= to_signed(0,32); mem_filters(21)(96) <= to_signed(0,32);
  mem_filters(21)(97) <= to_signed(0,32); mem_filters(21)(98) <= to_signed(0,32); mem_filters(21)(99) <= to_signed(0,32);
  mem_filters(21)(100) <= to_signed(0,32); mem_filters(21)(101) <= to_signed(0,32); mem_filters(21)(102) <= to_signed(0,32);
  mem_filters(21)(103) <= to_signed(0,32); mem_filters(21)(104) <= to_signed(0,32); mem_filters(21)(105) <= to_signed(0,32);
  mem_filters(21)(106) <= to_signed(0,32); mem_filters(21)(107) <= to_signed(0,32); mem_filters(21)(108) <= to_signed(0,32);
  mem_filters(21)(109) <= to_signed(0,32); mem_filters(21)(110) <= to_signed(0,32); mem_filters(21)(111) <= to_signed(0,32);
  mem_filters(21)(112) <= to_signed(0,32); mem_filters(21)(113) <= to_signed(0,32); mem_filters(21)(114) <= to_signed(0,32);
  mem_filters(21)(115) <= to_signed(0,32); mem_filters(21)(116) <= to_signed(0,32); mem_filters(21)(117) <= to_signed(0,32);
  mem_filters(21)(118) <= to_signed(0,32); mem_filters(21)(119) <= to_signed(0,32); mem_filters(21)(120) <= to_signed(0,32);
  mem_filters(21)(121) <= to_signed(0,32); mem_filters(21)(122) <= to_signed(0,32); mem_filters(21)(123) <= to_signed(0,32);
  mem_filters(21)(124) <= to_signed(0,32); mem_filters(21)(125) <= to_signed(0,32); mem_filters(21)(126) <= to_signed(0,32);
  mem_filters(21)(127) <= to_signed(0,32); mem_filters(21)(128) <= to_signed(0,32); mem_filters(21)(129) <= to_signed(0,32);
  mem_filters(21)(130) <= to_signed(0,32); mem_filters(21)(131) <= to_signed(0,32); mem_filters(21)(132) <= to_signed(0,32);
  mem_filters(21)(133) <= to_signed(0,32); mem_filters(21)(134) <= to_signed(0,32); mem_filters(21)(135) <= to_signed(0,32);
  mem_filters(21)(136) <= to_signed(0,32); mem_filters(21)(137) <= to_signed(0,32); mem_filters(21)(138) <= to_signed(0,32);
  mem_filters(21)(139) <= to_signed(0,32); mem_filters(21)(140) <= to_signed(0,32); mem_filters(21)(141) <= to_signed(0,32);
  mem_filters(21)(142) <= to_signed(0,32); mem_filters(21)(143) <= to_signed(0,32); mem_filters(21)(144) <= to_signed(0,32);
  mem_filters(21)(145) <= to_signed(0,32); mem_filters(21)(146) <= to_signed(0,32); mem_filters(21)(147) <= to_signed(0,32);
  mem_filters(21)(148) <= to_signed(0,32); mem_filters(21)(149) <= to_signed(0,32); mem_filters(21)(150) <= to_signed(0,32);
  mem_filters(21)(151) <= to_signed(0,32); mem_filters(21)(152) <= to_signed(0,32); mem_filters(21)(153) <= to_signed(0,32);
  mem_filters(21)(154) <= to_signed(0,32); mem_filters(21)(155) <= to_signed(0,32); mem_filters(21)(156) <= to_signed(0,32);
  mem_filters(21)(157) <= to_signed(0,32); mem_filters(21)(158) <= to_signed(0,32); mem_filters(21)(159) <= to_signed(0,32);
  mem_filters(21)(160) <= to_signed(0,32); mem_filters(21)(161) <= to_signed(0,32); mem_filters(21)(162) <= to_signed(0,32);
  mem_filters(21)(163) <= to_signed(0,32); mem_filters(21)(164) <= to_signed(0,32); mem_filters(21)(165) <= to_signed(0,32);
  mem_filters(21)(166) <= to_signed(0,32); mem_filters(21)(167) <= to_signed(0,32); mem_filters(21)(168) <= to_signed(0,32);
  mem_filters(21)(169) <= to_signed(0,32); mem_filters(21)(170) <= to_signed(0,32); mem_filters(21)(171) <= to_signed(0,32);
  mem_filters(21)(172) <= to_signed(0,32); mem_filters(21)(173) <= to_signed(0,32); mem_filters(21)(174) <= to_signed(0,32);
  mem_filters(21)(175) <= to_signed(0,32); mem_filters(21)(176) <= to_signed(0,32); mem_filters(21)(177) <= to_signed(0,32);
  mem_filters(21)(178) <= to_signed(0,32); mem_filters(21)(179) <= to_signed(0,32); mem_filters(21)(180) <= to_signed(0,32);
  mem_filters(21)(181) <= to_signed(0,32); mem_filters(21)(182) <= to_signed(0,32); mem_filters(21)(183) <= to_signed(0,32);
  mem_filters(21)(184) <= to_signed(0,32); mem_filters(21)(185) <= to_signed(0,32); mem_filters(21)(186) <= to_signed(0,32);
  mem_filters(21)(187) <= to_signed(0,32); mem_filters(21)(188) <= to_signed(0,32); mem_filters(21)(189) <= to_signed(0,32);
  mem_filters(21)(190) <= to_signed(0,32); mem_filters(21)(191) <= to_signed(0,32); mem_filters(21)(192) <= to_signed(0,32);
  mem_filters(21)(193) <= to_signed(0,32); mem_filters(21)(194) <= to_signed(0,32); mem_filters(21)(195) <= to_signed(0,32);
  mem_filters(21)(196) <= to_signed(0,32); mem_filters(21)(197) <= to_signed(0,32); mem_filters(21)(198) <= to_signed(0,32);
  mem_filters(21)(199) <= to_signed(0,32); mem_filters(21)(200) <= to_signed(0,32); mem_filters(21)(201) <= to_signed(0,32);
  mem_filters(21)(202) <= to_signed(0,32); mem_filters(21)(203) <= to_signed(0,32); mem_filters(21)(204) <= to_signed(0,32);
  mem_filters(21)(205) <= to_signed(0,32); mem_filters(21)(206) <= to_signed(0,32); mem_filters(21)(207) <= to_signed(0,32);
  mem_filters(21)(208) <= to_signed(0,32); mem_filters(21)(209) <= to_signed(0,32); mem_filters(21)(210) <= to_signed(0,32);
  mem_filters(21)(211) <= to_signed(0,32); mem_filters(21)(212) <= to_signed(0,32); mem_filters(21)(213) <= to_signed(0,32);
  mem_filters(21)(214) <= to_signed(0,32); mem_filters(21)(215) <= to_signed(0,32); mem_filters(21)(216) <= to_signed(0,32);
  mem_filters(21)(217) <= to_signed(0,32); mem_filters(21)(218) <= to_signed(0,32); mem_filters(21)(219) <= to_signed(0,32);
  mem_filters(21)(220) <= to_signed(0,32); mem_filters(21)(221) <= to_signed(0,32); mem_filters(21)(222) <= to_signed(0,32);
  mem_filters(21)(223) <= to_signed(0,32); mem_filters(21)(224) <= to_signed(0,32); mem_filters(21)(225) <= to_signed(0,32);
  mem_filters(21)(226) <= to_signed(0,32); mem_filters(21)(227) <= to_signed(0,32); mem_filters(21)(228) <= to_signed(0,32);
  mem_filters(21)(229) <= to_signed(0,32); mem_filters(21)(230) <= to_signed(0,32); mem_filters(21)(231) <= to_signed(0,32);
  mem_filters(21)(232) <= to_signed(0,32); mem_filters(21)(233) <= to_signed(0,32); mem_filters(21)(234) <= to_signed(0,32);
  mem_filters(21)(235) <= to_signed(0,32); mem_filters(21)(236) <= to_signed(0,32); mem_filters(21)(237) <= to_signed(0,32);
  mem_filters(21)(238) <= to_signed(0,32); mem_filters(21)(239) <= to_signed(0,32); mem_filters(21)(240) <= to_signed(0,32);
  mem_filters(21)(241) <= to_signed(0,32); mem_filters(21)(242) <= to_signed(0,32); mem_filters(21)(243) <= to_signed(0,32);
  mem_filters(21)(244) <= to_signed(0,32); mem_filters(21)(245) <= to_signed(0,32); mem_filters(21)(246) <= to_signed(0,32);
  mem_filters(21)(247) <= to_signed(0,32); mem_filters(21)(248) <= to_signed(0,32); mem_filters(21)(249) <= to_signed(0,32);
  mem_filters(21)(250) <= to_signed(0,32); mem_filters(21)(251) <= to_signed(0,32); mem_filters(21)(252) <= to_signed(0,32);
  mem_filters(21)(253) <= to_signed(0,32); mem_filters(21)(254) <= to_signed(0,32); mem_filters(21)(255) <= to_signed(0,32);
  
  --Filter 22
  mem_filters(22)(0) <= to_signed(0,32); mem_filters(22)(1) <= to_signed(0,32); mem_filters(22)(2) <= to_signed(0,32);
  mem_filters(22)(3) <= to_signed(0,32); mem_filters(22)(4) <= to_signed(0,32); mem_filters(22)(5) <= to_signed(0,32);
  mem_filters(22)(6) <= to_signed(0,32); mem_filters(22)(7) <= to_signed(0,32); mem_filters(22)(8) <= to_signed(0,32);
  mem_filters(22)(9) <= to_signed(0,32); mem_filters(22)(10) <= to_signed(0,32); mem_filters(22)(11) <= to_signed(0,32);
  mem_filters(22)(12) <= to_signed(0,32); mem_filters(22)(13) <= to_signed(0,32); mem_filters(22)(14) <= to_signed(0,32);
  mem_filters(22)(15) <= to_signed(0,32); mem_filters(22)(16) <= to_signed(0,32); mem_filters(22)(17) <= to_signed(0,32);
  mem_filters(22)(18) <= to_signed(0,32); mem_filters(22)(19) <= to_signed(0,32); mem_filters(22)(20) <= to_signed(0,32);
  mem_filters(22)(21) <= to_signed(0,32); mem_filters(22)(22) <= to_signed(0,32); mem_filters(22)(23) <= to_signed(0,32);
  mem_filters(22)(24) <= to_signed(0,32); mem_filters(22)(25) <= to_signed(0,32); mem_filters(22)(26) <= to_signed(0,32);
  mem_filters(22)(27) <= to_signed(0,32); mem_filters(22)(28) <= to_signed(0,32); mem_filters(22)(29) <= to_signed(0,32);
  mem_filters(22)(30) <= to_signed(0,32); mem_filters(22)(31) <= to_signed(0,32); mem_filters(22)(32) <= to_signed(0,32);
  mem_filters(22)(33) <= to_signed(0,32); mem_filters(22)(34) <= to_signed(0,32); mem_filters(22)(35) <= to_signed(0,32);
  mem_filters(22)(36) <= to_signed(0,32); mem_filters(22)(37) <= to_signed(0,32); mem_filters(22)(38) <= to_signed(0,32);
  mem_filters(22)(39) <= to_signed(0,32); mem_filters(22)(40) <= to_signed(0,32); mem_filters(22)(41) <= to_signed(0,32);
  mem_filters(22)(42) <= to_signed(0,32); mem_filters(22)(43) <= to_signed(0,32); mem_filters(22)(44) <= to_signed(0,32);
  mem_filters(22)(45) <= to_signed(0,32);
  mem_filters(22)(46) <= to_signed(0,32); mem_filters(22)(47) <= to_signed(0,32); mem_filters(22)(48) <= to_signed(0,32);
  mem_filters(22)(49) <= to_signed(0,32); mem_filters(22)(50) <= to_signed(0,32); mem_filters(22)(51) <= to_signed(0,32);
  mem_filters(22)(52) <= to_signed(0,32); mem_filters(22)(53) <= to_signed(0,32); mem_filters(22)(54) <= to_signed(0,32);
  mem_filters(22)(55) <= to_signed(0,32); mem_filters(22)(56) <= to_signed(0,32); mem_filters(22)(57) <= to_signed(0,32);
  mem_filters(22)(58) <= to_signed(0,32); mem_filters(22)(59) <= to_signed(0,32); mem_filters(22)(60) <= to_signed(0,32);
  mem_filters(22)(61) <= to_signed(0,32); mem_filters(22)(62) <= to_signed(0,32); mem_filters(22)(63) <= to_signed(0,32);
  mem_filters(22)(64) <= to_signed(0,32); mem_filters(22)(65) <= to_signed(0,32); mem_filters(22)(66) <= to_signed(0,32);
  mem_filters(22)(67) <= to_signed(0,32); mem_filters(22)(68) <= to_signed(0,32); mem_filters(22)(69) <= to_signed(0,32);
  mem_filters(22)(70) <= to_signed(0,32); mem_filters(22)(71) <= to_signed(0,32); mem_filters(22)(72) <= to_signed(0,32);
  mem_filters(22)(73) <= to_signed(0,32); mem_filters(22)(74) <= to_signed(0,32); mem_filters(22)(75) <= to_signed(0,32);
  mem_filters(22)(76) <= to_signed(0,32); mem_filters(22)(77) <= to_signed(0,32); mem_filters(22)(78) <= to_signed(0,32);
  mem_filters(22)(79) <= to_signed(0,32); mem_filters(22)(80) <= to_signed(0,32); mem_filters(22)(81) <= to_signed(0,32);
  mem_filters(22)(82) <= to_signed(0,32); mem_filters(22)(83) <= to_signed(0,32); mem_filters(22)(84) <= to_signed(0,32);
  mem_filters(22)(85) <= to_signed(0,32); mem_filters(22)(86) <= to_signed(0,32); mem_filters(22)(87) <= to_signed(0,32);
  mem_filters(22)(88) <= to_signed(0,32); mem_filters(22)(89) <= to_signed(0,32); mem_filters(22)(90) <= to_signed(0,32);
  mem_filters(22)(91) <= to_signed(0,32); mem_filters(22)(92) <= to_signed(0,32); mem_filters(22)(93) <= to_signed(0,32);
  mem_filters(22)(94) <= to_signed(0,32); mem_filters(22)(95) <= to_signed(0,32); mem_filters(22)(96) <= to_signed(0,32);
  mem_filters(22)(97) <= to_signed(0,32); mem_filters(22)(98) <= to_signed(0,32); mem_filters(22)(99) <= to_signed(0,32);
  mem_filters(22)(100) <= to_signed(0,32); mem_filters(22)(101) <= to_signed(0,32); mem_filters(22)(102) <= to_signed(0,32);
  mem_filters(22)(103) <= to_signed(0,32); mem_filters(22)(104) <= to_signed(0,32); mem_filters(22)(105) <= to_signed(0,32);
  mem_filters(22)(106) <= to_signed(0,32); mem_filters(22)(107) <= to_signed(0,32); mem_filters(22)(108) <= to_signed(0,32);
  mem_filters(22)(109) <= to_signed(0,32); mem_filters(22)(110) <= to_signed(0,32); mem_filters(22)(111) <= to_signed(0,32);
  mem_filters(22)(112) <= to_signed(0,32); mem_filters(22)(113) <= to_signed(0,32); mem_filters(22)(114) <= to_signed(0,32);
  mem_filters(22)(115) <= to_signed(0,32); mem_filters(22)(116) <= to_signed(0,32); mem_filters(22)(117) <= to_signed(0,32);
  mem_filters(22)(118) <= to_signed(0,32); mem_filters(22)(119) <= to_signed(0,32); mem_filters(22)(120) <= to_signed(0,32);
  mem_filters(22)(121) <= to_signed(0,32); mem_filters(22)(122) <= to_signed(0,32); mem_filters(22)(123) <= to_signed(0,32);
  mem_filters(22)(124) <= to_signed(0,32); mem_filters(22)(125) <= to_signed(0,32); mem_filters(22)(126) <= to_signed(0,32);
  mem_filters(22)(127) <= to_signed(0,32); mem_filters(22)(128) <= to_signed(0,32); mem_filters(22)(129) <= to_signed(0,32);
  mem_filters(22)(130) <= to_signed(0,32); mem_filters(22)(131) <= to_signed(0,32); mem_filters(22)(132) <= to_signed(0,32);
  mem_filters(22)(133) <= to_signed(0,32); mem_filters(22)(134) <= to_signed(0,32); mem_filters(22)(135) <= to_signed(0,32);
  mem_filters(22)(136) <= to_signed(0,32); mem_filters(22)(137) <= to_signed(0,32); mem_filters(22)(138) <= to_signed(0,32);
  mem_filters(22)(139) <= to_signed(0,32); mem_filters(22)(140) <= to_signed(0,32); mem_filters(22)(141) <= to_signed(0,32);
  mem_filters(22)(142) <= to_signed(0,32); mem_filters(22)(143) <= to_signed(0,32); mem_filters(22)(144) <= to_signed(0,32);
  mem_filters(22)(145) <= to_signed(0,32); mem_filters(22)(146) <= to_signed(0,32); mem_filters(22)(147) <= to_signed(0,32);
  mem_filters(22)(148) <= to_signed(0,32); mem_filters(22)(149) <= to_signed(0,32); mem_filters(22)(150) <= to_signed(0,32);
  mem_filters(22)(151) <= to_signed(0,32); mem_filters(22)(152) <= to_signed(0,32); mem_filters(22)(153) <= to_signed(0,32);
  mem_filters(22)(154) <= to_signed(0,32); mem_filters(22)(155) <= to_signed(0,32); mem_filters(22)(156) <= to_signed(0,32);
  mem_filters(22)(157) <= to_signed(0,32); mem_filters(22)(158) <= to_signed(0,32); mem_filters(22)(159) <= to_signed(0,32);
  mem_filters(22)(160) <= to_signed(0,32); mem_filters(22)(161) <= to_signed(0,32); mem_filters(22)(162) <= to_signed(0,32);
  mem_filters(22)(163) <= to_signed(0,32); mem_filters(22)(164) <= to_signed(0,32); mem_filters(22)(165) <= to_signed(0,32);
  mem_filters(22)(166) <= to_signed(0,32); mem_filters(22)(167) <= to_signed(0,32); mem_filters(22)(168) <= to_signed(0,32);
  mem_filters(22)(169) <= to_signed(0,32); mem_filters(22)(170) <= to_signed(0,32); mem_filters(22)(171) <= to_signed(0,32);
  mem_filters(22)(172) <= to_signed(0,32); mem_filters(22)(173) <= to_signed(0,32); mem_filters(22)(174) <= to_signed(0,32);
  mem_filters(22)(175) <= to_signed(0,32); mem_filters(22)(176) <= to_signed(0,32); mem_filters(22)(177) <= to_signed(0,32);
  mem_filters(22)(178) <= to_signed(0,32); mem_filters(22)(179) <= to_signed(0,32); mem_filters(22)(180) <= to_signed(0,32);
  mem_filters(22)(181) <= to_signed(0,32); mem_filters(22)(182) <= to_signed(0,32); mem_filters(22)(183) <= to_signed(0,32);
  mem_filters(22)(184) <= to_signed(0,32); mem_filters(22)(185) <= to_signed(0,32); mem_filters(22)(186) <= to_signed(0,32);
  mem_filters(22)(187) <= to_signed(0,32); mem_filters(22)(188) <= to_signed(0,32); mem_filters(22)(189) <= to_signed(0,32);
  mem_filters(22)(190) <= to_signed(0,32); mem_filters(22)(191) <= to_signed(0,32); mem_filters(22)(192) <= to_signed(0,32);
  mem_filters(22)(193) <= to_signed(0,32); mem_filters(22)(194) <= to_signed(0,32); mem_filters(22)(195) <= to_signed(0,32);
  mem_filters(22)(196) <= to_signed(0,32); mem_filters(22)(197) <= to_signed(0,32); mem_filters(22)(198) <= to_signed(0,32);
  mem_filters(22)(199) <= to_signed(0,32); mem_filters(22)(200) <= to_signed(0,32); mem_filters(22)(201) <= to_signed(0,32);
  mem_filters(22)(202) <= to_signed(0,32); mem_filters(22)(203) <= to_signed(0,32); mem_filters(22)(204) <= to_signed(0,32);
  mem_filters(22)(205) <= to_signed(0,32); mem_filters(22)(206) <= to_signed(0,32); mem_filters(22)(207) <= to_signed(0,32);
  mem_filters(22)(208) <= to_signed(0,32); mem_filters(22)(209) <= to_signed(0,32); mem_filters(22)(210) <= to_signed(0,32);
  mem_filters(22)(211) <= to_signed(0,32); mem_filters(22)(212) <= to_signed(0,32); mem_filters(22)(213) <= to_signed(0,32);
  mem_filters(22)(214) <= to_signed(0,32); mem_filters(22)(215) <= to_signed(0,32); mem_filters(22)(216) <= to_signed(0,32);
  mem_filters(22)(217) <= to_signed(0,32); mem_filters(22)(218) <= to_signed(0,32); mem_filters(22)(219) <= to_signed(0,32);
  mem_filters(22)(220) <= to_signed(0,32); mem_filters(22)(221) <= to_signed(0,32); mem_filters(22)(222) <= to_signed(0,32);
  mem_filters(22)(223) <= to_signed(0,32); mem_filters(22)(224) <= to_signed(0,32); mem_filters(22)(225) <= to_signed(0,32);
  mem_filters(22)(226) <= to_signed(0,32); mem_filters(22)(227) <= to_signed(0,32); mem_filters(22)(228) <= to_signed(0,32);
  mem_filters(22)(229) <= to_signed(0,32); mem_filters(22)(230) <= to_signed(0,32); mem_filters(22)(231) <= to_signed(0,32);
  mem_filters(22)(232) <= to_signed(0,32); mem_filters(22)(233) <= to_signed(0,32); mem_filters(22)(234) <= to_signed(0,32);
  mem_filters(22)(235) <= to_signed(0,32); mem_filters(22)(236) <= to_signed(0,32); mem_filters(22)(237) <= to_signed(0,32);
  mem_filters(22)(238) <= to_signed(0,32); mem_filters(22)(239) <= to_signed(0,32); mem_filters(22)(240) <= to_signed(0,32);
  mem_filters(22)(241) <= to_signed(0,32); mem_filters(22)(242) <= to_signed(0,32); mem_filters(22)(243) <= to_signed(0,32);
  mem_filters(22)(244) <= to_signed(0,32); mem_filters(22)(245) <= to_signed(0,32); mem_filters(22)(246) <= to_signed(0,32);
  mem_filters(22)(247) <= to_signed(0,32); mem_filters(22)(248) <= to_signed(0,32); mem_filters(22)(249) <= to_signed(0,32);
  mem_filters(22)(250) <= to_signed(0,32); mem_filters(22)(251) <= to_signed(0,32); mem_filters(22)(252) <= to_signed(0,32);
  mem_filters(22)(253) <= to_signed(0,32); mem_filters(22)(254) <= to_signed(0,32); mem_filters(22)(255) <= to_signed(0,32);
  
  --Filter 23
  mem_filters(23)(0) <= to_signed(0,32); mem_filters(23)(1) <= to_signed(0,32); mem_filters(23)(2) <= to_signed(0,32);
  mem_filters(23)(3) <= to_signed(0,32); mem_filters(23)(4) <= to_signed(0,32); mem_filters(23)(5) <= to_signed(0,32);
  mem_filters(23)(6) <= to_signed(0,32); mem_filters(23)(7) <= to_signed(0,32); mem_filters(23)(8) <= to_signed(0,32);
  mem_filters(23)(9) <= to_signed(0,32); mem_filters(23)(10) <= to_signed(0,32); mem_filters(23)(11) <= to_signed(0,32);
  mem_filters(23)(12) <= to_signed(0,32); mem_filters(23)(13) <= to_signed(0,32); mem_filters(23)(14) <= to_signed(0,32);
  mem_filters(23)(15) <= to_signed(0,32); mem_filters(23)(16) <= to_signed(0,32); mem_filters(23)(17) <= to_signed(0,32);
  mem_filters(23)(18) <= to_signed(0,32); mem_filters(23)(19) <= to_signed(0,32); mem_filters(23)(20) <= to_signed(0,32);
  mem_filters(23)(21) <= to_signed(0,32); mem_filters(23)(22) <= to_signed(0,32); mem_filters(23)(23) <= to_signed(0,32);
  mem_filters(23)(24) <= to_signed(0,32); mem_filters(23)(25) <= to_signed(0,32); mem_filters(23)(26) <= to_signed(0,32);
  mem_filters(23)(27) <= to_signed(0,32); mem_filters(23)(28) <= to_signed(0,32); mem_filters(23)(29) <= to_signed(0,32);
  mem_filters(23)(30) <= to_signed(0,32); mem_filters(23)(31) <= to_signed(0,32); mem_filters(23)(32) <= to_signed(0,32);
  mem_filters(23)(33) <= to_signed(0,32); mem_filters(23)(34) <= to_signed(0,32); mem_filters(23)(35) <= to_signed(0,32);
  mem_filters(23)(36) <= to_signed(0,32); mem_filters(23)(37) <= to_signed(0,32); mem_filters(23)(38) <= to_signed(0,32);
  mem_filters(23)(39) <= to_signed(0,32); mem_filters(23)(40) <= to_signed(0,32); mem_filters(23)(41) <= to_signed(0,32);
  mem_filters(23)(42) <= to_signed(0,32); mem_filters(23)(43) <= to_signed(0,32); mem_filters(23)(44) <= to_signed(0,32);
  mem_filters(23)(45) <= to_signed(0,32);
  mem_filters(23)(46) <= to_signed(0,32); mem_filters(23)(47) <= to_signed(0,32); mem_filters(23)(48) <= to_signed(0,32);
  mem_filters(23)(49) <= to_signed(0,32); mem_filters(23)(50) <= to_signed(0,32); mem_filters(23)(51) <= to_signed(0,32);
  mem_filters(23)(52) <= to_signed(0,32); mem_filters(23)(53) <= to_signed(0,32); mem_filters(23)(54) <= to_signed(0,32);
  mem_filters(23)(55) <= to_signed(0,32); mem_filters(23)(56) <= to_signed(0,32); mem_filters(23)(57) <= to_signed(0,32);
  mem_filters(23)(58) <= to_signed(0,32); mem_filters(23)(59) <= to_signed(0,32); mem_filters(23)(60) <= to_signed(0,32);
  mem_filters(23)(61) <= to_signed(0,32); mem_filters(23)(62) <= to_signed(0,32); mem_filters(23)(63) <= to_signed(0,32);
  mem_filters(23)(64) <= to_signed(0,32); mem_filters(23)(65) <= to_signed(0,32); mem_filters(23)(66) <= to_signed(0,32);
  mem_filters(23)(67) <= to_signed(0,32); mem_filters(23)(68) <= to_signed(0,32); mem_filters(23)(69) <= to_signed(0,32);
  mem_filters(23)(70) <= to_signed(0,32); mem_filters(23)(71) <= to_signed(0,32); mem_filters(23)(72) <= to_signed(0,32);
  mem_filters(23)(73) <= to_signed(0,32); mem_filters(23)(74) <= to_signed(0,32); mem_filters(23)(75) <= to_signed(0,32);
  mem_filters(23)(76) <= to_signed(0,32); mem_filters(23)(77) <= to_signed(0,32); mem_filters(23)(78) <= to_signed(0,32);
  mem_filters(23)(79) <= to_signed(0,32); mem_filters(23)(80) <= to_signed(0,32); mem_filters(23)(81) <= to_signed(0,32);
  mem_filters(23)(82) <= to_signed(0,32); mem_filters(23)(83) <= to_signed(0,32); mem_filters(23)(84) <= to_signed(0,32);
  mem_filters(23)(85) <= to_signed(0,32); mem_filters(23)(86) <= to_signed(0,32); mem_filters(23)(87) <= to_signed(0,32);
  mem_filters(23)(88) <= to_signed(0,32); mem_filters(23)(89) <= to_signed(0,32); mem_filters(23)(90) <= to_signed(0,32);
  mem_filters(23)(91) <= to_signed(0,32); mem_filters(23)(92) <= to_signed(0,32); mem_filters(23)(93) <= to_signed(0,32);
  mem_filters(23)(94) <= to_signed(0,32); mem_filters(23)(95) <= to_signed(0,32); mem_filters(23)(96) <= to_signed(0,32);
  mem_filters(23)(97) <= to_signed(0,32); mem_filters(23)(98) <= to_signed(0,32); mem_filters(23)(99) <= to_signed(0,32);
  mem_filters(23)(100) <= to_signed(0,32); mem_filters(23)(101) <= to_signed(0,32); mem_filters(23)(102) <= to_signed(0,32);
  mem_filters(23)(103) <= to_signed(0,32); mem_filters(23)(104) <= to_signed(0,32); mem_filters(23)(105) <= to_signed(0,32);
  mem_filters(23)(106) <= to_signed(0,32); mem_filters(23)(107) <= to_signed(0,32); mem_filters(23)(108) <= to_signed(0,32);
  mem_filters(23)(109) <= to_signed(0,32); mem_filters(23)(110) <= to_signed(0,32); mem_filters(23)(111) <= to_signed(0,32);
  mem_filters(23)(112) <= to_signed(0,32); mem_filters(23)(113) <= to_signed(0,32); mem_filters(23)(114) <= to_signed(0,32);
  mem_filters(23)(115) <= to_signed(0,32); mem_filters(23)(116) <= to_signed(0,32); mem_filters(23)(117) <= to_signed(0,32);
  mem_filters(23)(118) <= to_signed(0,32); mem_filters(23)(119) <= to_signed(0,32); mem_filters(23)(120) <= to_signed(0,32);
  mem_filters(23)(121) <= to_signed(0,32); mem_filters(23)(122) <= to_signed(0,32); mem_filters(23)(123) <= to_signed(0,32);
  mem_filters(23)(124) <= to_signed(0,32); mem_filters(23)(125) <= to_signed(0,32); mem_filters(23)(126) <= to_signed(0,32);
  mem_filters(23)(127) <= to_signed(0,32); mem_filters(23)(128) <= to_signed(0,32); mem_filters(23)(129) <= to_signed(0,32);
  mem_filters(23)(130) <= to_signed(0,32); mem_filters(23)(131) <= to_signed(0,32); mem_filters(23)(132) <= to_signed(0,32);
  mem_filters(23)(133) <= to_signed(0,32); mem_filters(23)(134) <= to_signed(0,32); mem_filters(23)(135) <= to_signed(0,32);
  mem_filters(23)(136) <= to_signed(0,32); mem_filters(23)(137) <= to_signed(0,32); mem_filters(23)(138) <= to_signed(0,32);
  mem_filters(23)(139) <= to_signed(0,32); mem_filters(23)(140) <= to_signed(0,32); mem_filters(23)(141) <= to_signed(0,32);
  mem_filters(23)(142) <= to_signed(0,32); mem_filters(23)(143) <= to_signed(0,32); mem_filters(23)(144) <= to_signed(0,32);
  mem_filters(23)(145) <= to_signed(0,32); mem_filters(23)(146) <= to_signed(0,32); mem_filters(23)(147) <= to_signed(0,32);
  mem_filters(23)(148) <= to_signed(0,32); mem_filters(23)(149) <= to_signed(0,32); mem_filters(23)(150) <= to_signed(0,32);
  mem_filters(23)(151) <= to_signed(0,32); mem_filters(23)(152) <= to_signed(0,32); mem_filters(23)(153) <= to_signed(0,32);
  mem_filters(23)(154) <= to_signed(0,32); mem_filters(23)(155) <= to_signed(0,32); mem_filters(23)(156) <= to_signed(0,32);
  mem_filters(23)(157) <= to_signed(0,32); mem_filters(23)(158) <= to_signed(0,32); mem_filters(23)(159) <= to_signed(0,32);
  mem_filters(23)(160) <= to_signed(0,32); mem_filters(23)(161) <= to_signed(0,32); mem_filters(23)(162) <= to_signed(0,32);
  mem_filters(23)(163) <= to_signed(0,32); mem_filters(23)(164) <= to_signed(0,32); mem_filters(23)(165) <= to_signed(0,32);
  mem_filters(23)(166) <= to_signed(0,32); mem_filters(23)(167) <= to_signed(0,32); mem_filters(23)(168) <= to_signed(0,32);
  mem_filters(23)(169) <= to_signed(0,32); mem_filters(23)(170) <= to_signed(0,32); mem_filters(23)(171) <= to_signed(0,32);
  mem_filters(23)(172) <= to_signed(0,32); mem_filters(23)(173) <= to_signed(0,32); mem_filters(23)(174) <= to_signed(0,32);
  mem_filters(23)(175) <= to_signed(0,32); mem_filters(23)(176) <= to_signed(0,32); mem_filters(23)(177) <= to_signed(0,32);
  mem_filters(23)(178) <= to_signed(0,32); mem_filters(23)(179) <= to_signed(0,32); mem_filters(23)(180) <= to_signed(0,32);
  mem_filters(23)(181) <= to_signed(0,32); mem_filters(23)(182) <= to_signed(0,32); mem_filters(23)(183) <= to_signed(0,32);
  mem_filters(23)(184) <= to_signed(0,32); mem_filters(23)(185) <= to_signed(0,32); mem_filters(23)(186) <= to_signed(0,32);
  mem_filters(23)(187) <= to_signed(0,32); mem_filters(23)(188) <= to_signed(0,32); mem_filters(23)(189) <= to_signed(0,32);
  mem_filters(23)(190) <= to_signed(0,32); mem_filters(23)(191) <= to_signed(0,32); mem_filters(23)(192) <= to_signed(0,32);
  mem_filters(23)(193) <= to_signed(0,32); mem_filters(23)(194) <= to_signed(0,32); mem_filters(23)(195) <= to_signed(0,32);
  mem_filters(23)(196) <= to_signed(0,32); mem_filters(23)(197) <= to_signed(0,32); mem_filters(23)(198) <= to_signed(0,32);
  mem_filters(23)(199) <= to_signed(0,32); mem_filters(23)(200) <= to_signed(0,32); mem_filters(23)(201) <= to_signed(0,32);
  mem_filters(23)(202) <= to_signed(0,32); mem_filters(23)(203) <= to_signed(0,32); mem_filters(23)(204) <= to_signed(0,32);
  mem_filters(23)(205) <= to_signed(0,32); mem_filters(23)(206) <= to_signed(0,32); mem_filters(23)(207) <= to_signed(0,32);
  mem_filters(23)(208) <= to_signed(0,32); mem_filters(23)(209) <= to_signed(0,32); mem_filters(23)(210) <= to_signed(0,32);
  mem_filters(23)(211) <= to_signed(0,32); mem_filters(23)(212) <= to_signed(0,32); mem_filters(23)(213) <= to_signed(0,32);
  mem_filters(23)(214) <= to_signed(0,32); mem_filters(23)(215) <= to_signed(0,32); mem_filters(23)(216) <= to_signed(0,32);
  mem_filters(23)(217) <= to_signed(0,32); mem_filters(23)(218) <= to_signed(0,32); mem_filters(23)(219) <= to_signed(0,32);
  mem_filters(23)(220) <= to_signed(0,32); mem_filters(23)(221) <= to_signed(0,32); mem_filters(23)(222) <= to_signed(0,32);
  mem_filters(23)(223) <= to_signed(0,32); mem_filters(23)(224) <= to_signed(0,32); mem_filters(23)(225) <= to_signed(0,32);
  mem_filters(23)(226) <= to_signed(0,32); mem_filters(23)(227) <= to_signed(0,32); mem_filters(23)(228) <= to_signed(0,32);
  mem_filters(23)(229) <= to_signed(0,32); mem_filters(23)(230) <= to_signed(0,32); mem_filters(23)(231) <= to_signed(0,32);
  mem_filters(23)(232) <= to_signed(0,32); mem_filters(23)(233) <= to_signed(0,32); mem_filters(23)(234) <= to_signed(0,32);
  mem_filters(23)(235) <= to_signed(0,32); mem_filters(23)(236) <= to_signed(0,32); mem_filters(23)(237) <= to_signed(0,32);
  mem_filters(23)(238) <= to_signed(0,32); mem_filters(23)(239) <= to_signed(0,32); mem_filters(23)(240) <= to_signed(0,32);
  mem_filters(23)(241) <= to_signed(0,32); mem_filters(23)(242) <= to_signed(0,32); mem_filters(23)(243) <= to_signed(0,32);
  mem_filters(23)(244) <= to_signed(0,32); mem_filters(23)(245) <= to_signed(0,32); mem_filters(23)(246) <= to_signed(0,32);
  mem_filters(23)(247) <= to_signed(0,32); mem_filters(23)(248) <= to_signed(0,32); mem_filters(23)(249) <= to_signed(0,32);
  mem_filters(23)(250) <= to_signed(0,32); mem_filters(23)(251) <= to_signed(0,32); mem_filters(23)(252) <= to_signed(0,32);
  mem_filters(23)(253) <= to_signed(0,32); mem_filters(23)(254) <= to_signed(0,32); mem_filters(23)(255) <= to_signed(0,32);
--end process;
end memery;