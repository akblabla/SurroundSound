library IEEE;
use IEEE.std_logic_1164.all;
use work.FilterTypes;

entity FilterInterpolator is
	port(test : in std_logic);
end entity FilterInterpolator;

architecture default of FilterInterpolator is
begin
end default;