library IEEE;
use IEEE.std_logic_1164.all;
use work.FilterTypes;

entity SurroundSound is
	port(test : in std_logic);
end entity SurroundSound;

architecture default of SurroundSound is
begin
end default;